`timescale 1 ns / 1 ps 

module fmm_reduce_kernel_greedy_potential_reduce_with_debug_Pipeline_VITIS_LOOP_135_110 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        new_col_3,
        mul_ln132,
        M_e_address0,
        M_e_ce0,
        M_e_we0,
        M_e_d0,
        M_e_address1,
        M_e_ce1,
        M_e_q1,
        mul_ln133,
        mul_ln144,
        icmp_ln133,
        cmp34_i_i
);

parameter    ap_ST_fsm_pp0_stage0 = 3'd1;
parameter    ap_ST_fsm_pp0_stage1 = 3'd2;
parameter    ap_ST_fsm_pp0_stage2 = 3'd4;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [31:0] new_col_3;
input  [16:0] mul_ln132;
output  [16:0] M_e_address0;
output   M_e_ce0;
output   M_e_we0;
output  [31:0] M_e_d0;
output  [16:0] M_e_address1;
output   M_e_ce1;
input  [31:0] M_e_q1;
input  [16:0] mul_ln133;
input  [16:0] mul_ln144;
input  [0:0] icmp_ln133;
input  [0:0] cmp34_i_i;

reg ap_idle;

(* fsm_encoding = "none" *) reg   [2:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
reg    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_idle_pp0;
wire    ap_CS_fsm_pp0_stage2;
wire    ap_block_pp0_stage2_subdone;
reg    ap_enable_reg_pp0_iter0_reg;
reg   [0:0] icmp_ln135_reg_242;
reg    ap_condition_exit_pp0_iter0_stage2;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln135_fu_131_p2;
wire   [16:0] trunc_ln137_fu_143_p1;
reg   [16:0] trunc_ln137_reg_246;
reg   [16:0] M_e_addr_5_reg_252;
reg   [16:0] M_e_addr_7_reg_258;
wire    ap_CS_fsm_pp0_stage1;
wire    ap_block_pp0_stage1_11001;
reg   [16:0] M_e_addr_reg_264;
reg   [16:0] M_e_addr_reg_264_pp0_iter1_reg;
reg  signed [31:0] e1_reg_269;
reg  signed [31:0] e1_reg_269_pp0_iter1_reg;
wire   [0:0] grp_fu_113_p2;
reg   [0:0] icmp_ln138_reg_276;
reg   [0:0] icmp_ln140_reg_280;
wire    ap_block_pp0_stage2_11001;
wire   [0:0] and_ln141_fu_186_p2;
reg   [0:0] and_ln141_reg_284;
wire   [0:0] or_ln141_fu_191_p2;
reg   [0:0] or_ln141_reg_288;
wire   [0:0] icmp_ln141_1_fu_209_p2;
reg   [0:0] icmp_ln141_1_reg_292;
wire   [63:0] zext_ln137_fu_153_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln139_fu_167_p1;
wire    ap_block_pp0_stage1;
wire   [63:0] zext_ln144_fu_176_p1;
reg   [30:0] c_2_fu_40;
wire   [30:0] add_ln135_fu_137_p2;
wire    ap_loop_init;
reg   [30:0] ap_sig_allocacmp_c;
reg    M_e_ce1_local;
reg   [16:0] M_e_address1_local;
reg    M_e_we0_local;
reg   [31:0] M_e_d0_local;
reg    M_e_ce0_local;
reg   [16:0] M_e_address0_local;
reg    ap_predicate_pred177_state5;
reg    ap_predicate_pred177_state6;
wire    ap_block_pp0_stage2;
wire  signed [31:0] grp_fu_113_p0;
wire   [31:0] zext_ln135_fu_127_p1;
wire   [16:0] add_ln137_fu_147_p2;
wire   [16:0] add_ln139_fu_163_p2;
wire   [16:0] add_ln144_fu_172_p2;
wire  signed [31:0] icmp_ln141_fu_181_p1;
wire   [0:0] icmp_ln141_fu_181_p2;
wire  signed [31:0] sext_ln141_fu_196_p0;
wire  signed [32:0] sext_ln141_fu_196_p1;
wire  signed [32:0] sext_ln141_1_fu_206_p1;
wire   [32:0] sub_ln141_fu_200_p2;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg   [2:0] ap_NS_fsm;
wire    ap_block_pp0_stage0_subdone;
reg    ap_idle_pp0_1to1;
wire    ap_block_pp0_stage1_subdone;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ready_sig;
wire    ap_done_sig;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 3'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter0_reg = 1'b0;
#0 c_2_fu_40 = 31'd0;
#0 ap_done_reg = 1'b0;
end

fmm_reduce_kernel_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready_sig),
    .ap_done(ap_done_sig),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter0_stage2),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter0_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
            ap_enable_reg_pp0_iter0_reg <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter0_stage2)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            ap_enable_reg_pp0_iter1 <= ap_enable_reg_pp0_iter0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if (((icmp_ln135_fu_131_p2 == 1'd1) & (ap_enable_reg_pp0_iter0 == 1'b1))) begin
            c_2_fu_40 <= add_ln135_fu_137_p2;
        end else if ((ap_loop_init == 1'b1)) begin
            c_2_fu_40 <= 31'd0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        M_e_addr_5_reg_252 <= zext_ln137_fu_153_p1;
        ap_predicate_pred177_state5 <= (((icmp_ln141_1_reg_292 == 1'd1) & (or_ln141_reg_288 == 1'd0) & (icmp_ln140_reg_280 == 1'd0) & (icmp_ln138_reg_276 == 1'd0)) | ((1'd1 == and_ln141_reg_284) & (or_ln141_reg_288 == 1'd1) & (icmp_ln140_reg_280 == 1'd0) & (icmp_ln138_reg_276 == 1'd0)));
        icmp_ln135_reg_242 <= icmp_ln135_fu_131_p2;
        trunc_ln137_reg_246 <= trunc_ln137_fu_143_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        M_e_addr_7_reg_258 <= zext_ln139_fu_167_p1;
        M_e_addr_reg_264 <= zext_ln144_fu_176_p1;
        M_e_addr_reg_264_pp0_iter1_reg <= M_e_addr_reg_264;
        ap_predicate_pred177_state6 <= (((icmp_ln141_1_reg_292 == 1'd1) & (or_ln141_reg_288 == 1'd0) & (icmp_ln140_reg_280 == 1'd0) & (icmp_ln138_reg_276 == 1'd0)) | ((1'd1 == and_ln141_reg_284) & (or_ln141_reg_288 == 1'd1) & (icmp_ln140_reg_280 == 1'd0) & (icmp_ln138_reg_276 == 1'd0)));
        e1_reg_269_pp0_iter1_reg <= e1_reg_269;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        and_ln141_reg_284 <= and_ln141_fu_186_p2;
        icmp_ln141_1_reg_292 <= icmp_ln141_1_fu_209_p2;
        or_ln141_reg_288 <= or_ln141_fu_191_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0_reg == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        e1_reg_269 <= M_e_q1;
        icmp_ln138_reg_276 <= grp_fu_113_p2;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0_reg == 1'b1) & (1'b0 == ap_block_pp0_stage2_11001) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        icmp_ln140_reg_280 <= grp_fu_113_p2;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
        if (((1'b0 == ap_block_pp0_stage2) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
            M_e_address0_local = M_e_addr_reg_264_pp0_iter1_reg;
        end else if (((1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
            M_e_address0_local = M_e_addr_7_reg_258;
        end else if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            M_e_address0_local = M_e_addr_5_reg_252;
        end else begin
            M_e_address0_local = 'bx;
        end
    end else begin
        M_e_address0_local = 'bx;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0_reg == 1'b1) & (1'b0 == ap_block_pp0_stage1) & (1'b1 == ap_CS_fsm_pp0_stage1))) begin
        M_e_address1_local = zext_ln139_fu_167_p1;
    end else if (((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        M_e_address1_local = zext_ln137_fu_153_p1;
    end else begin
        M_e_address1_local = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2)))) begin
        M_e_ce0_local = 1'b1;
    end else begin
        M_e_ce0_local = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)) | ((ap_enable_reg_pp0_iter0_reg == 1'b1) & (1'b0 == ap_block_pp0_stage1_11001) & (1'b1 == ap_CS_fsm_pp0_stage1)))) begin
        M_e_ce1_local = 1'b1;
    end else begin
        M_e_ce1_local = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage2) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        M_e_d0_local = e1_reg_269_pp0_iter1_reg;
    end else if ((((1'b0 == ap_block_pp0_stage1) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1)) | ((1'b0 == ap_block_pp0_stage0) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0)))) begin
        M_e_d0_local = 32'd0;
    end else begin
        M_e_d0_local = 'bx;
    end
end

always @ (*) begin
    if ((((1'b0 == ap_block_pp0_stage1_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage1) & (ap_predicate_pred177_state5 == 1'b1)) | ((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (((icmp_ln141_1_reg_292 == 1'd1) & (or_ln141_reg_288 == 1'd0) & (icmp_ln140_reg_280 == 1'd0) & (icmp_ln138_reg_276 == 1'd0)) | ((1'd1 == and_ln141_reg_284) & (or_ln141_reg_288 == 1'd1) & (icmp_ln140_reg_280 == 1'd0) & (icmp_ln138_reg_276 == 1'd0)))) | ((1'b0 == ap_block_pp0_stage2_11001) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage2) & (ap_predicate_pred177_state6 == 1'b1)))) begin
        M_e_we0_local = 1'b1;
    end else begin
        M_e_we0_local = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln135_reg_242 == 1'd0) & (ap_enable_reg_pp0_iter0_reg == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        ap_condition_exit_pp0_iter0_stage2 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter0_stage2 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_pp0_stage0)) begin
        ap_enable_reg_pp0_iter0 = ap_start_int;
    end else begin
        ap_enable_reg_pp0_iter0 = ap_enable_reg_pp0_iter0_reg;
    end
end

always @ (*) begin
    if (((ap_start_int == 1'b0) & (ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if ((ap_enable_reg_pp0_iter1 == 1'b0)) begin
        ap_idle_pp0_1to1 = 1'b1;
    end else begin
        ap_idle_pp0_1to1 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0_reg == 1'b1) & (1'b0 == ap_block_pp0_stage2_subdone) & (1'b1 == ap_CS_fsm_pp0_stage2))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
        ap_sig_allocacmp_c = 31'd0;
    end else begin
        ap_sig_allocacmp_c = c_2_fu_40;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            if ((~((ap_start_int == 1'b0) & (ap_idle_pp0_1to1 == 1'b1)) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end
        end
        ap_ST_fsm_pp0_stage1 : begin
            if ((1'b0 == ap_block_pp0_stage1_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage1;
            end
        end
        ap_ST_fsm_pp0_stage2 : begin
            if ((1'b0 == ap_block_pp0_stage2_subdone)) begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage0;
            end else begin
                ap_NS_fsm = ap_ST_fsm_pp0_stage2;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign M_e_address0 = M_e_address0_local;

assign M_e_address1 = M_e_address1_local;

assign M_e_ce0 = M_e_ce0_local;

assign M_e_ce1 = M_e_ce1_local;

assign M_e_d0 = M_e_d0_local;

assign M_e_we0 = M_e_we0_local;

assign add_ln135_fu_137_p2 = (ap_sig_allocacmp_c + 31'd1);

assign add_ln137_fu_147_p2 = (mul_ln132 + trunc_ln137_fu_143_p1);

assign add_ln139_fu_163_p2 = (mul_ln133 + trunc_ln137_reg_246);

assign add_ln144_fu_172_p2 = (mul_ln144 + trunc_ln137_reg_246);

assign and_ln141_fu_186_p2 = (icmp_ln141_fu_181_p2 & icmp_ln133);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_pp0_stage1 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_pp0_stage2 = ap_CS_fsm[32'd2];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage1_subdone = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage2_subdone = ~(1'b1 == 1'b1);

assign ap_done = ap_done_sig;

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter0_stage2;

assign ap_ready = ap_ready_sig;

assign grp_fu_113_p0 = M_e_q1;

assign grp_fu_113_p2 = ((grp_fu_113_p0 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln135_fu_131_p2 = (($signed(zext_ln135_fu_127_p1) < $signed(new_col_3)) ? 1'b1 : 1'b0);

assign icmp_ln141_1_fu_209_p2 = ((sext_ln141_1_fu_206_p1 == sub_ln141_fu_200_p2) ? 1'b1 : 1'b0);

assign icmp_ln141_fu_181_p1 = M_e_q1;

assign icmp_ln141_fu_181_p2 = ((e1_reg_269 == icmp_ln141_fu_181_p1) ? 1'b1 : 1'b0);

assign or_ln141_fu_191_p2 = (cmp34_i_i | and_ln141_fu_186_p2);

assign sext_ln141_1_fu_206_p1 = e1_reg_269;

assign sext_ln141_fu_196_p0 = M_e_q1;

assign sext_ln141_fu_196_p1 = sext_ln141_fu_196_p0;

assign sub_ln141_fu_200_p2 = ($signed(33'd0) - $signed(sext_ln141_fu_196_p1));

assign trunc_ln137_fu_143_p1 = ap_sig_allocacmp_c[16:0];

assign zext_ln135_fu_127_p1 = ap_sig_allocacmp_c;

assign zext_ln137_fu_153_p1 = add_ln137_fu_147_p2;

assign zext_ln139_fu_167_p1 = add_ln139_fu_163_p2;

assign zext_ln144_fu_176_p1 = add_ln144_fu_172_p2;

endmodule //fmm_reduce_kernel_greedy_potential_reduce_with_debug_Pipeline_VITIS_LOOP_135_110
