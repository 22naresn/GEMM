`timescale 1 ns / 1 ps 

module fmm_reduce_kernel_load_matrix_from_dram_safe (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_gmem_0_AWVALID,
        m_axi_gmem_0_AWREADY,
        m_axi_gmem_0_AWADDR,
        m_axi_gmem_0_AWID,
        m_axi_gmem_0_AWLEN,
        m_axi_gmem_0_AWSIZE,
        m_axi_gmem_0_AWBURST,
        m_axi_gmem_0_AWLOCK,
        m_axi_gmem_0_AWCACHE,
        m_axi_gmem_0_AWPROT,
        m_axi_gmem_0_AWQOS,
        m_axi_gmem_0_AWREGION,
        m_axi_gmem_0_AWUSER,
        m_axi_gmem_0_WVALID,
        m_axi_gmem_0_WREADY,
        m_axi_gmem_0_WDATA,
        m_axi_gmem_0_WSTRB,
        m_axi_gmem_0_WLAST,
        m_axi_gmem_0_WID,
        m_axi_gmem_0_WUSER,
        m_axi_gmem_0_ARVALID,
        m_axi_gmem_0_ARREADY,
        m_axi_gmem_0_ARADDR,
        m_axi_gmem_0_ARID,
        m_axi_gmem_0_ARLEN,
        m_axi_gmem_0_ARSIZE,
        m_axi_gmem_0_ARBURST,
        m_axi_gmem_0_ARLOCK,
        m_axi_gmem_0_ARCACHE,
        m_axi_gmem_0_ARPROT,
        m_axi_gmem_0_ARQOS,
        m_axi_gmem_0_ARREGION,
        m_axi_gmem_0_ARUSER,
        m_axi_gmem_0_RVALID,
        m_axi_gmem_0_RREADY,
        m_axi_gmem_0_RDATA,
        m_axi_gmem_0_RLAST,
        m_axi_gmem_0_RID,
        m_axi_gmem_0_RFIFONUM,
        m_axi_gmem_0_RUSER,
        m_axi_gmem_0_RRESP,
        m_axi_gmem_0_BVALID,
        m_axi_gmem_0_BREADY,
        m_axi_gmem_0_BRESP,
        m_axi_gmem_0_BID,
        m_axi_gmem_0_BUSER,
        A_dram,
        rows,
        cols,
        t_capacity,
        M_e_address0,
        M_e_ce0,
        M_e_we0,
        M_e_d0,
        M_rows,
        M_rows_ap_vld,
        M_cols,
        M_cols_ap_vld,
        M_t,
        M_t_ap_vld,
        M_t_capacity,
        M_t_capacity_ap_vld
);

parameter    ap_ST_fsm_state1 = 4'd1;
parameter    ap_ST_fsm_state2 = 4'd2;
parameter    ap_ST_fsm_state3 = 4'd4;
parameter    ap_ST_fsm_state4 = 4'd8;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_gmem_0_AWVALID;
input   m_axi_gmem_0_AWREADY;
output  [63:0] m_axi_gmem_0_AWADDR;
output  [0:0] m_axi_gmem_0_AWID;
output  [31:0] m_axi_gmem_0_AWLEN;
output  [2:0] m_axi_gmem_0_AWSIZE;
output  [1:0] m_axi_gmem_0_AWBURST;
output  [1:0] m_axi_gmem_0_AWLOCK;
output  [3:0] m_axi_gmem_0_AWCACHE;
output  [2:0] m_axi_gmem_0_AWPROT;
output  [3:0] m_axi_gmem_0_AWQOS;
output  [3:0] m_axi_gmem_0_AWREGION;
output  [0:0] m_axi_gmem_0_AWUSER;
output   m_axi_gmem_0_WVALID;
input   m_axi_gmem_0_WREADY;
output  [31:0] m_axi_gmem_0_WDATA;
output  [3:0] m_axi_gmem_0_WSTRB;
output   m_axi_gmem_0_WLAST;
output  [0:0] m_axi_gmem_0_WID;
output  [0:0] m_axi_gmem_0_WUSER;
output   m_axi_gmem_0_ARVALID;
input   m_axi_gmem_0_ARREADY;
output  [63:0] m_axi_gmem_0_ARADDR;
output  [0:0] m_axi_gmem_0_ARID;
output  [31:0] m_axi_gmem_0_ARLEN;
output  [2:0] m_axi_gmem_0_ARSIZE;
output  [1:0] m_axi_gmem_0_ARBURST;
output  [1:0] m_axi_gmem_0_ARLOCK;
output  [3:0] m_axi_gmem_0_ARCACHE;
output  [2:0] m_axi_gmem_0_ARPROT;
output  [3:0] m_axi_gmem_0_ARQOS;
output  [3:0] m_axi_gmem_0_ARREGION;
output  [0:0] m_axi_gmem_0_ARUSER;
input   m_axi_gmem_0_RVALID;
output   m_axi_gmem_0_RREADY;
input  [31:0] m_axi_gmem_0_RDATA;
input   m_axi_gmem_0_RLAST;
input  [0:0] m_axi_gmem_0_RID;
input  [8:0] m_axi_gmem_0_RFIFONUM;
input  [0:0] m_axi_gmem_0_RUSER;
input  [1:0] m_axi_gmem_0_RRESP;
input   m_axi_gmem_0_BVALID;
output   m_axi_gmem_0_BREADY;
input  [1:0] m_axi_gmem_0_BRESP;
input  [0:0] m_axi_gmem_0_BID;
input  [0:0] m_axi_gmem_0_BUSER;
input  [63:0] A_dram;
input  [31:0] rows;
input  [31:0] cols;
input  [31:0] t_capacity;
output  [16:0] M_e_address0;
output   M_e_ce0;
output   M_e_we0;
output  [31:0] M_e_d0;
output  [31:0] M_rows;
output   M_rows_ap_vld;
output  [31:0] M_cols;
output   M_cols_ap_vld;
output  [31:0] M_t;
output   M_t_ap_vld;
output  [31:0] M_t_capacity;
output   M_t_capacity_ap_vld;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg[16:0] M_e_address0;
reg M_e_ce0;
reg M_e_we0;
reg[31:0] M_e_d0;
reg M_rows_ap_vld;
reg M_cols_ap_vld;
reg M_t_ap_vld;
reg M_t_capacity_ap_vld;

(* fsm_encoding = "none" *) reg   [3:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
wire   [30:0] smax_fu_121_p3;
reg   [30:0] smax_reg_169;
wire   [30:0] smax2_fu_135_p3;
reg   [30:0] smax2_reg_174;
wire   [61:0] mul_ln58_fu_91_p2;
reg   [61:0] mul_ln58_reg_179;
wire    ap_CS_fsm_state2;
wire    ap_CS_fsm_state3;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_start;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_done;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_idle;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_ready;
wire   [16:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_address0;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_ce0;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_we0;
wire   [31:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_d0;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_start;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_done;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_idle;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_ready;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWVALID;
wire   [63:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWADDR;
wire   [0:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWID;
wire   [31:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWLEN;
wire   [2:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWSIZE;
wire   [1:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWBURST;
wire   [1:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWLOCK;
wire   [3:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWCACHE;
wire   [2:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWPROT;
wire   [3:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWQOS;
wire   [3:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWREGION;
wire   [0:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWUSER;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WVALID;
wire   [31:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WDATA;
wire   [3:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WSTRB;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WLAST;
wire   [0:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WID;
wire   [0:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WUSER;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARVALID;
wire   [63:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARADDR;
wire   [0:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARID;
wire   [31:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARLEN;
wire   [2:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARSIZE;
wire   [1:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARBURST;
wire   [1:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARLOCK;
wire   [3:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARCACHE;
wire   [2:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARPROT;
wire   [3:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARQOS;
wire   [3:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARREGION;
wire   [0:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARUSER;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_RREADY;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_BREADY;
wire   [16:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_address0;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_ce0;
wire    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_we0;
wire   [31:0] grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_d0;
reg    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_start_reg;
reg    grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_start_reg;
wire    ap_CS_fsm_state4;
wire   [30:0] mul_ln58_fu_91_p0;
wire   [30:0] mul_ln58_fu_91_p1;
wire   [0:0] empty_41_fu_115_p2;
wire   [30:0] empty_40_fu_99_p1;
wire   [0:0] empty_42_fu_129_p2;
wire   [30:0] empty_fu_95_p1;
reg   [3:0] ap_NS_fsm;
reg    ap_ST_fsm_state1_blk;
reg    ap_ST_fsm_state2_blk;
wire    ap_ST_fsm_state3_blk;
reg    ap_ST_fsm_state4_blk;
wire   [61:0] mul_ln58_fu_91_p00;
wire   [61:0] mul_ln58_fu_91_p10;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 4'd1;
#0 grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_start_reg = 1'b0;
#0 grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_start_reg = 1'b0;
end

fmm_reduce_kernel_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2 grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_start),
    .ap_done(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_done),
    .ap_idle(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_idle),
    .ap_ready(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_ready),
    .M_e_address0(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_address0),
    .M_e_ce0(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_ce0),
    .M_e_we0(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_we0),
    .M_e_d0(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_d0)
);

fmm_reduce_kernel_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4 grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_start),
    .ap_done(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_done),
    .ap_idle(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_idle),
    .ap_ready(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_ready),
    .m_axi_gmem_0_AWVALID(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWVALID),
    .m_axi_gmem_0_AWREADY(1'b0),
    .m_axi_gmem_0_AWADDR(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWADDR),
    .m_axi_gmem_0_AWID(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWID),
    .m_axi_gmem_0_AWLEN(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWLEN),
    .m_axi_gmem_0_AWSIZE(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWSIZE),
    .m_axi_gmem_0_AWBURST(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWBURST),
    .m_axi_gmem_0_AWLOCK(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWLOCK),
    .m_axi_gmem_0_AWCACHE(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWCACHE),
    .m_axi_gmem_0_AWPROT(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWPROT),
    .m_axi_gmem_0_AWQOS(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWQOS),
    .m_axi_gmem_0_AWREGION(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWREGION),
    .m_axi_gmem_0_AWUSER(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_AWUSER),
    .m_axi_gmem_0_WVALID(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WVALID),
    .m_axi_gmem_0_WREADY(1'b0),
    .m_axi_gmem_0_WDATA(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WDATA),
    .m_axi_gmem_0_WSTRB(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WSTRB),
    .m_axi_gmem_0_WLAST(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WLAST),
    .m_axi_gmem_0_WID(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WID),
    .m_axi_gmem_0_WUSER(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_WUSER),
    .m_axi_gmem_0_ARVALID(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARVALID),
    .m_axi_gmem_0_ARREADY(m_axi_gmem_0_ARREADY),
    .m_axi_gmem_0_ARADDR(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARADDR),
    .m_axi_gmem_0_ARID(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARID),
    .m_axi_gmem_0_ARLEN(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARLEN),
    .m_axi_gmem_0_ARSIZE(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARSIZE),
    .m_axi_gmem_0_ARBURST(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARBURST),
    .m_axi_gmem_0_ARLOCK(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARLOCK),
    .m_axi_gmem_0_ARCACHE(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARCACHE),
    .m_axi_gmem_0_ARPROT(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARPROT),
    .m_axi_gmem_0_ARQOS(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARQOS),
    .m_axi_gmem_0_ARREGION(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARREGION),
    .m_axi_gmem_0_ARUSER(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARUSER),
    .m_axi_gmem_0_RVALID(m_axi_gmem_0_RVALID),
    .m_axi_gmem_0_RREADY(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_RREADY),
    .m_axi_gmem_0_RDATA(m_axi_gmem_0_RDATA),
    .m_axi_gmem_0_RLAST(m_axi_gmem_0_RLAST),
    .m_axi_gmem_0_RID(m_axi_gmem_0_RID),
    .m_axi_gmem_0_RFIFONUM(m_axi_gmem_0_RFIFONUM),
    .m_axi_gmem_0_RUSER(m_axi_gmem_0_RUSER),
    .m_axi_gmem_0_RRESP(m_axi_gmem_0_RRESP),
    .m_axi_gmem_0_BVALID(1'b0),
    .m_axi_gmem_0_BREADY(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_BREADY),
    .m_axi_gmem_0_BRESP(2'd0),
    .m_axi_gmem_0_BID(1'd0),
    .m_axi_gmem_0_BUSER(1'd0),
    .cols(cols),
    .mul_ln58(mul_ln58_reg_179),
    .A_dram(A_dram),
    .sext_ln58(cols),
    .M_e_address0(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_address0),
    .M_e_ce0(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_ce0),
    .M_e_we0(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_we0),
    .M_e_d0(grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_d0)
);

fmm_reduce_kernel_mul_31ns_31ns_62_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 31 ),
    .din1_WIDTH( 31 ),
    .dout_WIDTH( 62 ))
mul_31ns_31ns_62_1_1_U28(
    .din0(mul_ln58_fu_91_p0),
    .din1(mul_ln58_fu_91_p1),
    .dout(mul_ln58_fu_91_p2)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_start_reg <= 1'b0;
    end else begin
        if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
            grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_start_reg <= 1'b1;
        end else if ((grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_ready == 1'b1)) begin
            grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state3)) begin
            grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_start_reg <= 1'b1;
        end else if ((grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_ready == 1'b1)) begin
            grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        mul_ln58_reg_179 <= mul_ln58_fu_91_p2;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b1 == ap_CS_fsm_state1)) begin
        smax2_reg_174 <= smax2_fu_135_p3;
        smax_reg_169 <= smax_fu_121_p3;
    end
end

always @ (*) begin
    if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        M_cols_ap_vld = 1'b1;
    end else begin
        M_cols_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        M_e_address0 = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_address0;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        M_e_address0 = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_address0;
    end else begin
        M_e_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        M_e_ce0 = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_ce0;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        M_e_ce0 = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_ce0;
    end else begin
        M_e_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        M_e_d0 = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_d0;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        M_e_d0 = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_d0;
    end else begin
        M_e_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state4)) begin
        M_e_we0 = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_M_e_we0;
    end else if ((1'b1 == ap_CS_fsm_state2)) begin
        M_e_we0 = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_M_e_we0;
    end else begin
        M_e_we0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
        M_rows_ap_vld = 1'b1;
    end else begin
        M_rows_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_done == 1'b1))) begin
        M_t_ap_vld = 1'b1;
    end else begin
        M_t_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_done == 1'b1))) begin
        M_t_capacity_ap_vld = 1'b1;
    end else begin
        M_t_capacity_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if ((ap_start == 1'b0)) begin
        ap_ST_fsm_state1_blk = 1'b1;
    end else begin
        ap_ST_fsm_state1_blk = 1'b0;
    end
end

always @ (*) begin
    if ((grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_done == 1'b0)) begin
        ap_ST_fsm_state2_blk = 1'b1;
    end else begin
        ap_ST_fsm_state2_blk = 1'b0;
    end
end

assign ap_ST_fsm_state3_blk = 1'b0;

always @ (*) begin
    if ((grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_done == 1'b0)) begin
        ap_ST_fsm_state4_blk = 1'b1;
    end else begin
        ap_ST_fsm_state4_blk = 1'b0;
    end
end

always @ (*) begin
    if ((((1'b1 == ap_CS_fsm_state4) & (grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_done == 1'b1)) | ((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1)))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = 1'b0;
    end
end

always @ (*) begin
    if (((ap_start == 1'b0) & (1'b1 == ap_CS_fsm_state1))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state4) & (grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_done == 1'b1))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((ap_start == 1'b1) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((1'b1 == ap_CS_fsm_state2) & (grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_done == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
        end
        ap_ST_fsm_state3 : begin
            ap_NS_fsm = ap_ST_fsm_state4;
        end
        ap_ST_fsm_state4 : begin
            if (((1'b1 == ap_CS_fsm_state4) & (grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_done == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign M_cols = cols;

assign M_rows = rows;

assign M_t = 32'd0;

assign M_t_capacity = t_capacity;

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state4 = ap_CS_fsm[32'd3];

assign empty_40_fu_99_p1 = rows[30:0];

assign empty_41_fu_115_p2 = (($signed(rows) > $signed(32'd0)) ? 1'b1 : 1'b0);

assign empty_42_fu_129_p2 = (($signed(cols) > $signed(32'd0)) ? 1'b1 : 1'b0);

assign empty_fu_95_p1 = cols[30:0];

assign grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_start = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2_fu_72_ap_start_reg;

assign grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_start = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_ap_start_reg;

assign m_axi_gmem_0_ARADDR = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARADDR;

assign m_axi_gmem_0_ARBURST = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARBURST;

assign m_axi_gmem_0_ARCACHE = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARCACHE;

assign m_axi_gmem_0_ARID = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARID;

assign m_axi_gmem_0_ARLEN = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARLEN;

assign m_axi_gmem_0_ARLOCK = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARLOCK;

assign m_axi_gmem_0_ARPROT = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARPROT;

assign m_axi_gmem_0_ARQOS = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARQOS;

assign m_axi_gmem_0_ARREGION = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARREGION;

assign m_axi_gmem_0_ARSIZE = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARSIZE;

assign m_axi_gmem_0_ARUSER = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARUSER;

assign m_axi_gmem_0_ARVALID = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_ARVALID;

assign m_axi_gmem_0_AWADDR = 64'd0;

assign m_axi_gmem_0_AWBURST = 2'd0;

assign m_axi_gmem_0_AWCACHE = 4'd0;

assign m_axi_gmem_0_AWID = 1'd0;

assign m_axi_gmem_0_AWLEN = 32'd0;

assign m_axi_gmem_0_AWLOCK = 2'd0;

assign m_axi_gmem_0_AWPROT = 3'd0;

assign m_axi_gmem_0_AWQOS = 4'd0;

assign m_axi_gmem_0_AWREGION = 4'd0;

assign m_axi_gmem_0_AWSIZE = 3'd0;

assign m_axi_gmem_0_AWUSER = 1'd0;

assign m_axi_gmem_0_AWVALID = 1'b0;

assign m_axi_gmem_0_BREADY = 1'b0;

assign m_axi_gmem_0_RREADY = grp_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4_fu_78_m_axi_gmem_0_RREADY;

assign m_axi_gmem_0_WDATA = 32'd0;

assign m_axi_gmem_0_WID = 1'd0;

assign m_axi_gmem_0_WLAST = 1'b0;

assign m_axi_gmem_0_WSTRB = 4'd0;

assign m_axi_gmem_0_WUSER = 1'd0;

assign m_axi_gmem_0_WVALID = 1'b0;

assign mul_ln58_fu_91_p0 = mul_ln58_fu_91_p00;

assign mul_ln58_fu_91_p00 = smax_reg_169;

assign mul_ln58_fu_91_p1 = mul_ln58_fu_91_p10;

assign mul_ln58_fu_91_p10 = smax2_reg_174;

assign smax2_fu_135_p3 = ((empty_42_fu_129_p2[0:0] == 1'b1) ? empty_fu_95_p1 : 31'd0);

assign smax_fu_121_p3 = ((empty_41_fu_115_p2[0:0] == 1'b1) ? empty_40_fu_99_p1 : 31'd0);

endmodule //fmm_reduce_kernel_load_matrix_from_dram_safe
