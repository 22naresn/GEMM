`timescale 1 ns / 1 ps 

module fmm_reduce_kernel_Block_entry_proc (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_continue,
        ap_idle,
        ap_ready,
        p_read,
        p_read1,
        m_axi_gmem_0_AWVALID,
        m_axi_gmem_0_AWREADY,
        m_axi_gmem_0_AWADDR,
        m_axi_gmem_0_AWID,
        m_axi_gmem_0_AWLEN,
        m_axi_gmem_0_AWSIZE,
        m_axi_gmem_0_AWBURST,
        m_axi_gmem_0_AWLOCK,
        m_axi_gmem_0_AWCACHE,
        m_axi_gmem_0_AWPROT,
        m_axi_gmem_0_AWQOS,
        m_axi_gmem_0_AWREGION,
        m_axi_gmem_0_AWUSER,
        m_axi_gmem_0_WVALID,
        m_axi_gmem_0_WREADY,
        m_axi_gmem_0_WDATA,
        m_axi_gmem_0_WSTRB,
        m_axi_gmem_0_WLAST,
        m_axi_gmem_0_WID,
        m_axi_gmem_0_WUSER,
        m_axi_gmem_0_ARVALID,
        m_axi_gmem_0_ARREADY,
        m_axi_gmem_0_ARADDR,
        m_axi_gmem_0_ARID,
        m_axi_gmem_0_ARLEN,
        m_axi_gmem_0_ARSIZE,
        m_axi_gmem_0_ARBURST,
        m_axi_gmem_0_ARLOCK,
        m_axi_gmem_0_ARCACHE,
        m_axi_gmem_0_ARPROT,
        m_axi_gmem_0_ARQOS,
        m_axi_gmem_0_ARREGION,
        m_axi_gmem_0_ARUSER,
        m_axi_gmem_0_RVALID,
        m_axi_gmem_0_RREADY,
        m_axi_gmem_0_RDATA,
        m_axi_gmem_0_RLAST,
        m_axi_gmem_0_RID,
        m_axi_gmem_0_RFIFONUM,
        m_axi_gmem_0_RUSER,
        m_axi_gmem_0_RRESP,
        m_axi_gmem_0_BVALID,
        m_axi_gmem_0_BREADY,
        m_axi_gmem_0_BRESP,
        m_axi_gmem_0_BID,
        m_axi_gmem_0_BUSER,
        A_dram_dout,
        A_dram_empty_n,
        A_dram_read,
        A_dram_num_data_valid,
        A_dram_fifo_cap,
        rows_dout,
        rows_empty_n,
        rows_read,
        rows_num_data_valid,
        rows_fifo_cap,
        cols_dout,
        cols_empty_n,
        cols_read,
        cols_num_data_valid,
        cols_fifo_cap,
        t_capacity_dout,
        t_capacity_empty_n,
        t_capacity_read,
        t_capacity_num_data_valid,
        t_capacity_fifo_cap,
        k1_dout,
        k1_empty_n,
        k1_read,
        k1_num_data_valid,
        k1_fifo_cap,
        k2_dout,
        k2_empty_n,
        k2_read,
        k2_num_data_valid,
        k2_fifo_cap,
        m_axi_gmem2_0_AWVALID,
        m_axi_gmem2_0_AWREADY,
        m_axi_gmem2_0_AWADDR,
        m_axi_gmem2_0_AWID,
        m_axi_gmem2_0_AWLEN,
        m_axi_gmem2_0_AWSIZE,
        m_axi_gmem2_0_AWBURST,
        m_axi_gmem2_0_AWLOCK,
        m_axi_gmem2_0_AWCACHE,
        m_axi_gmem2_0_AWPROT,
        m_axi_gmem2_0_AWQOS,
        m_axi_gmem2_0_AWREGION,
        m_axi_gmem2_0_AWUSER,
        m_axi_gmem2_0_WVALID,
        m_axi_gmem2_0_WREADY,
        m_axi_gmem2_0_WDATA,
        m_axi_gmem2_0_WSTRB,
        m_axi_gmem2_0_WLAST,
        m_axi_gmem2_0_WID,
        m_axi_gmem2_0_WUSER,
        m_axi_gmem2_0_ARVALID,
        m_axi_gmem2_0_ARREADY,
        m_axi_gmem2_0_ARADDR,
        m_axi_gmem2_0_ARID,
        m_axi_gmem2_0_ARLEN,
        m_axi_gmem2_0_ARSIZE,
        m_axi_gmem2_0_ARBURST,
        m_axi_gmem2_0_ARLOCK,
        m_axi_gmem2_0_ARCACHE,
        m_axi_gmem2_0_ARPROT,
        m_axi_gmem2_0_ARQOS,
        m_axi_gmem2_0_ARREGION,
        m_axi_gmem2_0_ARUSER,
        m_axi_gmem2_0_RVALID,
        m_axi_gmem2_0_RREADY,
        m_axi_gmem2_0_RDATA,
        m_axi_gmem2_0_RLAST,
        m_axi_gmem2_0_RID,
        m_axi_gmem2_0_RFIFONUM,
        m_axi_gmem2_0_RUSER,
        m_axi_gmem2_0_RRESP,
        m_axi_gmem2_0_BVALID,
        m_axi_gmem2_0_BREADY,
        m_axi_gmem2_0_BRESP,
        m_axi_gmem2_0_BID,
        m_axi_gmem2_0_BUSER,
        debug_dram_dout,
        debug_dram_empty_n,
        debug_dram_read,
        debug_dram_num_data_valid,
        debug_dram_fifo_cap,
        debug_capacity_dout,
        debug_capacity_empty_n,
        debug_capacity_read,
        debug_capacity_num_data_valid,
        debug_capacity_fifo_cap
);

parameter    ap_ST_fsm_state1 = 13'd1;
parameter    ap_ST_fsm_state2 = 13'd2;
parameter    ap_ST_fsm_state3 = 13'd4;
parameter    ap_ST_fsm_state4 = 13'd8;
parameter    ap_ST_fsm_state5 = 13'd16;
parameter    ap_ST_fsm_state6 = 13'd32;
parameter    ap_ST_fsm_state7 = 13'd64;
parameter    ap_ST_fsm_state8 = 13'd128;
parameter    ap_ST_fsm_state9 = 13'd256;
parameter    ap_ST_fsm_state10 = 13'd512;
parameter    ap_ST_fsm_state11 = 13'd1024;
parameter    ap_ST_fsm_state12 = 13'd2048;
parameter    ap_ST_fsm_state13 = 13'd4096;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
input   ap_continue;
output   ap_idle;
output   ap_ready;
input  [0:0] p_read;
input  [0:0] p_read1;
output   m_axi_gmem_0_AWVALID;
input   m_axi_gmem_0_AWREADY;
output  [63:0] m_axi_gmem_0_AWADDR;
output  [0:0] m_axi_gmem_0_AWID;
output  [31:0] m_axi_gmem_0_AWLEN;
output  [2:0] m_axi_gmem_0_AWSIZE;
output  [1:0] m_axi_gmem_0_AWBURST;
output  [1:0] m_axi_gmem_0_AWLOCK;
output  [3:0] m_axi_gmem_0_AWCACHE;
output  [2:0] m_axi_gmem_0_AWPROT;
output  [3:0] m_axi_gmem_0_AWQOS;
output  [3:0] m_axi_gmem_0_AWREGION;
output  [0:0] m_axi_gmem_0_AWUSER;
output   m_axi_gmem_0_WVALID;
input   m_axi_gmem_0_WREADY;
output  [31:0] m_axi_gmem_0_WDATA;
output  [3:0] m_axi_gmem_0_WSTRB;
output   m_axi_gmem_0_WLAST;
output  [0:0] m_axi_gmem_0_WID;
output  [0:0] m_axi_gmem_0_WUSER;
output   m_axi_gmem_0_ARVALID;
input   m_axi_gmem_0_ARREADY;
output  [63:0] m_axi_gmem_0_ARADDR;
output  [0:0] m_axi_gmem_0_ARID;
output  [31:0] m_axi_gmem_0_ARLEN;
output  [2:0] m_axi_gmem_0_ARSIZE;
output  [1:0] m_axi_gmem_0_ARBURST;
output  [1:0] m_axi_gmem_0_ARLOCK;
output  [3:0] m_axi_gmem_0_ARCACHE;
output  [2:0] m_axi_gmem_0_ARPROT;
output  [3:0] m_axi_gmem_0_ARQOS;
output  [3:0] m_axi_gmem_0_ARREGION;
output  [0:0] m_axi_gmem_0_ARUSER;
input   m_axi_gmem_0_RVALID;
output   m_axi_gmem_0_RREADY;
input  [31:0] m_axi_gmem_0_RDATA;
input   m_axi_gmem_0_RLAST;
input  [0:0] m_axi_gmem_0_RID;
input  [8:0] m_axi_gmem_0_RFIFONUM;
input  [0:0] m_axi_gmem_0_RUSER;
input  [1:0] m_axi_gmem_0_RRESP;
input   m_axi_gmem_0_BVALID;
output   m_axi_gmem_0_BREADY;
input  [1:0] m_axi_gmem_0_BRESP;
input  [0:0] m_axi_gmem_0_BID;
input  [0:0] m_axi_gmem_0_BUSER;
input  [63:0] A_dram_dout;
input   A_dram_empty_n;
output   A_dram_read;
input  [2:0] A_dram_num_data_valid;
input  [2:0] A_dram_fifo_cap;
input  [31:0] rows_dout;
input   rows_empty_n;
output   rows_read;
input  [2:0] rows_num_data_valid;
input  [2:0] rows_fifo_cap;
input  [31:0] cols_dout;
input   cols_empty_n;
output   cols_read;
input  [2:0] cols_num_data_valid;
input  [2:0] cols_fifo_cap;
input  [31:0] t_capacity_dout;
input   t_capacity_empty_n;
output   t_capacity_read;
input  [2:0] t_capacity_num_data_valid;
input  [2:0] t_capacity_fifo_cap;
input  [31:0] k1_dout;
input   k1_empty_n;
output   k1_read;
input  [2:0] k1_num_data_valid;
input  [2:0] k1_fifo_cap;
input  [31:0] k2_dout;
input   k2_empty_n;
output   k2_read;
input  [2:0] k2_num_data_valid;
input  [2:0] k2_fifo_cap;
output   m_axi_gmem2_0_AWVALID;
input   m_axi_gmem2_0_AWREADY;
output  [63:0] m_axi_gmem2_0_AWADDR;
output  [0:0] m_axi_gmem2_0_AWID;
output  [31:0] m_axi_gmem2_0_AWLEN;
output  [2:0] m_axi_gmem2_0_AWSIZE;
output  [1:0] m_axi_gmem2_0_AWBURST;
output  [1:0] m_axi_gmem2_0_AWLOCK;
output  [3:0] m_axi_gmem2_0_AWCACHE;
output  [2:0] m_axi_gmem2_0_AWPROT;
output  [3:0] m_axi_gmem2_0_AWQOS;
output  [3:0] m_axi_gmem2_0_AWREGION;
output  [0:0] m_axi_gmem2_0_AWUSER;
output   m_axi_gmem2_0_WVALID;
input   m_axi_gmem2_0_WREADY;
output  [31:0] m_axi_gmem2_0_WDATA;
output  [3:0] m_axi_gmem2_0_WSTRB;
output   m_axi_gmem2_0_WLAST;
output  [0:0] m_axi_gmem2_0_WID;
output  [0:0] m_axi_gmem2_0_WUSER;
output   m_axi_gmem2_0_ARVALID;
input   m_axi_gmem2_0_ARREADY;
output  [63:0] m_axi_gmem2_0_ARADDR;
output  [0:0] m_axi_gmem2_0_ARID;
output  [31:0] m_axi_gmem2_0_ARLEN;
output  [2:0] m_axi_gmem2_0_ARSIZE;
output  [1:0] m_axi_gmem2_0_ARBURST;
output  [1:0] m_axi_gmem2_0_ARLOCK;
output  [3:0] m_axi_gmem2_0_ARCACHE;
output  [2:0] m_axi_gmem2_0_ARPROT;
output  [3:0] m_axi_gmem2_0_ARQOS;
output  [3:0] m_axi_gmem2_0_ARREGION;
output  [0:0] m_axi_gmem2_0_ARUSER;
input   m_axi_gmem2_0_RVALID;
output   m_axi_gmem2_0_RREADY;
input  [31:0] m_axi_gmem2_0_RDATA;
input   m_axi_gmem2_0_RLAST;
input  [0:0] m_axi_gmem2_0_RID;
input  [8:0] m_axi_gmem2_0_RFIFONUM;
input  [0:0] m_axi_gmem2_0_RUSER;
input  [1:0] m_axi_gmem2_0_RRESP;
input   m_axi_gmem2_0_BVALID;
output   m_axi_gmem2_0_BREADY;
input  [1:0] m_axi_gmem2_0_BRESP;
input  [0:0] m_axi_gmem2_0_BID;
input  [0:0] m_axi_gmem2_0_BUSER;
input  [63:0] debug_dram_dout;
input   debug_dram_empty_n;
output   debug_dram_read;
input  [2:0] debug_dram_num_data_valid;
input  [2:0] debug_dram_fifo_cap;
input  [31:0] debug_capacity_dout;
input   debug_capacity_empty_n;
output   debug_capacity_read;
input  [2:0] debug_capacity_num_data_valid;
input  [2:0] debug_capacity_fifo_cap;

reg ap_done;
reg ap_idle;
reg ap_ready;
reg m_axi_gmem_0_AWVALID;
reg m_axi_gmem_0_WVALID;
reg m_axi_gmem_0_ARVALID;
reg m_axi_gmem_0_RREADY;
reg m_axi_gmem_0_BREADY;
reg A_dram_read;
reg rows_read;
reg cols_read;
reg t_capacity_read;
reg k1_read;
reg k2_read;
reg m_axi_gmem2_0_AWVALID;
reg[63:0] m_axi_gmem2_0_AWADDR;
reg[0:0] m_axi_gmem2_0_AWID;
reg[31:0] m_axi_gmem2_0_AWLEN;
reg[2:0] m_axi_gmem2_0_AWSIZE;
reg[1:0] m_axi_gmem2_0_AWBURST;
reg[1:0] m_axi_gmem2_0_AWLOCK;
reg[3:0] m_axi_gmem2_0_AWCACHE;
reg[2:0] m_axi_gmem2_0_AWPROT;
reg[3:0] m_axi_gmem2_0_AWQOS;
reg[3:0] m_axi_gmem2_0_AWREGION;
reg[0:0] m_axi_gmem2_0_AWUSER;
reg m_axi_gmem2_0_WVALID;
reg[31:0] m_axi_gmem2_0_WDATA;
reg[3:0] m_axi_gmem2_0_WSTRB;
reg m_axi_gmem2_0_WLAST;
reg[0:0] m_axi_gmem2_0_WID;
reg[0:0] m_axi_gmem2_0_WUSER;
reg m_axi_gmem2_0_BREADY;
reg debug_dram_read;
reg debug_capacity_read;

reg    ap_done_reg;
(* fsm_encoding = "none" *) reg   [12:0] ap_CS_fsm;
wire    ap_CS_fsm_state1;
reg   [31:0] M_rows;
reg   [31:0] M_cols;
reg   [31:0] M_t;
reg   [31:0] M_t_capacity;
reg   [16:0] M_e_address0;
reg    M_e_ce0;
reg    M_e_we0;
reg   [31:0] M_e_d0;
wire   [31:0] M_e_q0;
reg    M_e_ce1;
reg    M_e_we1;
wire   [31:0] M_e_q1;
reg    A_dram_blk_n;
reg    rows_blk_n;
reg    cols_blk_n;
reg    t_capacity_blk_n;
reg    k1_blk_n;
reg    k2_blk_n;
reg    gmem2_blk_n_AW;
wire    ap_CS_fsm_state2;
reg    gmem2_blk_n_W;
wire    ap_CS_fsm_state3;
reg    gmem2_blk_n_B;
wire    ap_CS_fsm_state8;
reg   [0:0] and_ln307_reg_317;
reg   [0:0] icmp_ln308_reg_321;
reg    debug_dram_blk_n;
reg    debug_capacity_blk_n;
reg   [0:0] p_read_2_reg_270;
reg    ap_block_state1;
reg   [31:0] debug_capacity_read_reg_275;
reg   [63:0] debug_dram_read_reg_280;
reg   [31:0] k2_read_reg_286;
reg   [31:0] k1_read_reg_291;
reg   [31:0] t_capacity_read_reg_296;
reg   [31:0] cols_read_reg_301;
reg   [31:0] rows_read_reg_306;
reg   [63:0] A_dram_read_reg_311;
wire   [0:0] and_ln307_fu_231_p2;
wire   [0:0] icmp_ln308_fu_237_p2;
wire   [31:0] select_ln309_fu_243_p3;
reg   [31:0] select_ln309_reg_325;
wire    grp_load_matrix_from_dram_safe_fu_174_ap_start;
wire    grp_load_matrix_from_dram_safe_fu_174_ap_done;
wire    grp_load_matrix_from_dram_safe_fu_174_ap_idle;
wire    grp_load_matrix_from_dram_safe_fu_174_ap_ready;
wire    grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWVALID;
wire   [63:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWADDR;
wire   [0:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWID;
wire   [31:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWLEN;
wire   [2:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWSIZE;
wire   [1:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWBURST;
wire   [1:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWLOCK;
wire   [3:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWCACHE;
wire   [2:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWPROT;
wire   [3:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWQOS;
wire   [3:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWREGION;
wire   [0:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWUSER;
wire    grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WVALID;
wire   [31:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WDATA;
wire   [3:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WSTRB;
wire    grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WLAST;
wire   [0:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WID;
wire   [0:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WUSER;
wire    grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARVALID;
wire   [63:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARADDR;
wire   [0:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARID;
wire   [31:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARLEN;
wire   [2:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARSIZE;
wire   [1:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARBURST;
wire   [1:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARLOCK;
wire   [3:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARCACHE;
wire   [2:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARPROT;
wire   [3:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARQOS;
wire   [3:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARREGION;
wire   [0:0] grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARUSER;
wire    grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_RREADY;
wire    grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_BREADY;
wire   [16:0] grp_load_matrix_from_dram_safe_fu_174_M_e_address0;
wire    grp_load_matrix_from_dram_safe_fu_174_M_e_ce0;
wire    grp_load_matrix_from_dram_safe_fu_174_M_e_we0;
wire   [31:0] grp_load_matrix_from_dram_safe_fu_174_M_e_d0;
wire   [31:0] grp_load_matrix_from_dram_safe_fu_174_M_rows;
wire    grp_load_matrix_from_dram_safe_fu_174_M_rows_ap_vld;
wire   [31:0] grp_load_matrix_from_dram_safe_fu_174_M_cols;
wire    grp_load_matrix_from_dram_safe_fu_174_M_cols_ap_vld;
wire   [31:0] grp_load_matrix_from_dram_safe_fu_174_M_t;
wire    grp_load_matrix_from_dram_safe_fu_174_M_t_ap_vld;
wire   [31:0] grp_load_matrix_from_dram_safe_fu_174_M_t_capacity;
wire    grp_load_matrix_from_dram_safe_fu_174_M_t_capacity_ap_vld;
wire    grp_greedy_potential_reduce_with_debug_fu_198_ap_start;
wire    grp_greedy_potential_reduce_with_debug_fu_198_ap_done;
wire    grp_greedy_potential_reduce_with_debug_fu_198_ap_idle;
wire    grp_greedy_potential_reduce_with_debug_fu_198_ap_ready;
wire    grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWVALID;
wire   [63:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWADDR;
wire   [0:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWID;
wire   [31:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWLEN;
wire   [2:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWSIZE;
wire   [1:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWBURST;
wire   [1:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWLOCK;
wire   [3:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWCACHE;
wire   [2:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWPROT;
wire   [3:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWQOS;
wire   [3:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWREGION;
wire   [0:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWUSER;
wire    grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WVALID;
wire   [31:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WDATA;
wire   [3:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WSTRB;
wire    grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WLAST;
wire   [0:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WID;
wire   [0:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WUSER;
wire    grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARVALID;
wire   [63:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARADDR;
wire   [0:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARID;
wire   [31:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARLEN;
wire   [2:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARSIZE;
wire   [1:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARBURST;
wire   [1:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARLOCK;
wire   [3:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARCACHE;
wire   [2:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARPROT;
wire   [3:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARQOS;
wire   [3:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARREGION;
wire   [0:0] grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARUSER;
wire    grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_RREADY;
wire    grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_BREADY;
wire   [16:0] grp_greedy_potential_reduce_with_debug_fu_198_M_e_address0;
wire    grp_greedy_potential_reduce_with_debug_fu_198_M_e_ce0;
wire    grp_greedy_potential_reduce_with_debug_fu_198_M_e_we0;
wire   [31:0] grp_greedy_potential_reduce_with_debug_fu_198_M_e_d0;
wire   [16:0] grp_greedy_potential_reduce_with_debug_fu_198_M_e_address1;
wire    grp_greedy_potential_reduce_with_debug_fu_198_M_e_ce1;
wire    grp_greedy_potential_reduce_with_debug_fu_198_M_e_we1;
wire   [31:0] grp_greedy_potential_reduce_with_debug_fu_198_M_e_d1;
wire   [31:0] grp_greedy_potential_reduce_with_debug_fu_198_M_t_o;
wire    grp_greedy_potential_reduce_with_debug_fu_198_M_t_o_ap_vld;
wire    grp_store_matrix_to_dram_safe_fu_218_ap_start;
wire    grp_store_matrix_to_dram_safe_fu_218_ap_done;
wire    grp_store_matrix_to_dram_safe_fu_218_ap_idle;
wire    grp_store_matrix_to_dram_safe_fu_218_ap_ready;
wire    grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWVALID;
wire   [63:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWADDR;
wire   [0:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWID;
wire   [31:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWLEN;
wire   [2:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWSIZE;
wire   [1:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWBURST;
wire   [1:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWLOCK;
wire   [3:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWCACHE;
wire   [2:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWPROT;
wire   [3:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWQOS;
wire   [3:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWREGION;
wire   [0:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWUSER;
wire    grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WVALID;
wire   [31:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WDATA;
wire   [3:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WSTRB;
wire    grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WLAST;
wire   [0:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WID;
wire   [0:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WUSER;
wire    grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARVALID;
wire   [63:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARADDR;
wire   [0:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARID;
wire   [31:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARLEN;
wire   [2:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARSIZE;
wire   [1:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARBURST;
wire   [1:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARLOCK;
wire   [3:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARCACHE;
wire   [2:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARPROT;
wire   [3:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARQOS;
wire   [3:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARREGION;
wire   [0:0] grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARUSER;
wire    grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_RREADY;
wire    grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_BREADY;
wire   [16:0] grp_store_matrix_to_dram_safe_fu_218_M_e_address0;
wire    grp_store_matrix_to_dram_safe_fu_218_M_e_ce0;
reg    grp_load_matrix_from_dram_safe_fu_174_ap_start_reg;
reg    ap_block_state1_ignore_call0;
wire    ap_CS_fsm_state9;
reg    grp_greedy_potential_reduce_with_debug_fu_198_ap_start_reg;
wire    ap_CS_fsm_state10;
wire    ap_CS_fsm_state11;
reg    grp_store_matrix_to_dram_safe_fu_218_ap_start_reg;
wire    ap_CS_fsm_state12;
wire    ap_CS_fsm_state13;
wire  signed [63:0] sext_ln309_fu_259_p1;
reg    ap_predicate_op49_writeresp_state8;
reg    ap_block_state8;
wire   [61:0] trunc_ln_fu_250_p4;
reg   [12:0] ap_NS_fsm;
reg    ap_ST_fsm_state1_blk;
reg    ap_ST_fsm_state2_blk;
reg    ap_ST_fsm_state3_blk;
wire    ap_ST_fsm_state4_blk;
wire    ap_ST_fsm_state5_blk;
wire    ap_ST_fsm_state6_blk;
wire    ap_ST_fsm_state7_blk;
reg    ap_ST_fsm_state8_blk;
reg    ap_ST_fsm_state9_blk;
wire    ap_ST_fsm_state10_blk;
reg    ap_ST_fsm_state11_blk;
wire    ap_ST_fsm_state12_blk;
reg    ap_ST_fsm_state13_blk;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_done_reg = 1'b0;
#0 ap_CS_fsm = 13'd1;
#0 M_rows = 32'd0;
#0 M_cols = 32'd0;
#0 M_t = 32'd0;
#0 M_t_capacity = 32'd0;
#0 grp_load_matrix_from_dram_safe_fu_174_ap_start_reg = 1'b0;
#0 grp_greedy_potential_reduce_with_debug_fu_198_ap_start_reg = 1'b0;
#0 grp_store_matrix_to_dram_safe_fu_218_ap_start_reg = 1'b0;
end

fmm_reduce_kernel_Block_entry_proc_M_e_RAM_AUTO_1R1W #(
    .DataWidth( 32 ),
    .AddressRange( 102400 ),
    .AddressWidth( 17 ))
M_e_U(
    .clk(ap_clk),
    .reset(ap_rst),
    .address0(M_e_address0),
    .ce0(M_e_ce0),
    .we0(M_e_we0),
    .d0(M_e_d0),
    .q0(M_e_q0),
    .address1(grp_greedy_potential_reduce_with_debug_fu_198_M_e_address1),
    .ce1(M_e_ce1),
    .we1(M_e_we1),
    .d1(grp_greedy_potential_reduce_with_debug_fu_198_M_e_d1),
    .q1(M_e_q1)
);

fmm_reduce_kernel_load_matrix_from_dram_safe grp_load_matrix_from_dram_safe_fu_174(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_load_matrix_from_dram_safe_fu_174_ap_start),
    .ap_done(grp_load_matrix_from_dram_safe_fu_174_ap_done),
    .ap_idle(grp_load_matrix_from_dram_safe_fu_174_ap_idle),
    .ap_ready(grp_load_matrix_from_dram_safe_fu_174_ap_ready),
    .m_axi_gmem_0_AWVALID(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWVALID),
    .m_axi_gmem_0_AWREADY(1'b0),
    .m_axi_gmem_0_AWADDR(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWADDR),
    .m_axi_gmem_0_AWID(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWID),
    .m_axi_gmem_0_AWLEN(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWLEN),
    .m_axi_gmem_0_AWSIZE(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWSIZE),
    .m_axi_gmem_0_AWBURST(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWBURST),
    .m_axi_gmem_0_AWLOCK(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWLOCK),
    .m_axi_gmem_0_AWCACHE(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWCACHE),
    .m_axi_gmem_0_AWPROT(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWPROT),
    .m_axi_gmem_0_AWQOS(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWQOS),
    .m_axi_gmem_0_AWREGION(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWREGION),
    .m_axi_gmem_0_AWUSER(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_AWUSER),
    .m_axi_gmem_0_WVALID(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WVALID),
    .m_axi_gmem_0_WREADY(1'b0),
    .m_axi_gmem_0_WDATA(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WDATA),
    .m_axi_gmem_0_WSTRB(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WSTRB),
    .m_axi_gmem_0_WLAST(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WLAST),
    .m_axi_gmem_0_WID(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WID),
    .m_axi_gmem_0_WUSER(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_WUSER),
    .m_axi_gmem_0_ARVALID(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARVALID),
    .m_axi_gmem_0_ARREADY(m_axi_gmem_0_ARREADY),
    .m_axi_gmem_0_ARADDR(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARADDR),
    .m_axi_gmem_0_ARID(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARID),
    .m_axi_gmem_0_ARLEN(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARLEN),
    .m_axi_gmem_0_ARSIZE(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARSIZE),
    .m_axi_gmem_0_ARBURST(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARBURST),
    .m_axi_gmem_0_ARLOCK(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARLOCK),
    .m_axi_gmem_0_ARCACHE(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARCACHE),
    .m_axi_gmem_0_ARPROT(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARPROT),
    .m_axi_gmem_0_ARQOS(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARQOS),
    .m_axi_gmem_0_ARREGION(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARREGION),
    .m_axi_gmem_0_ARUSER(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARUSER),
    .m_axi_gmem_0_RVALID(m_axi_gmem_0_RVALID),
    .m_axi_gmem_0_RREADY(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_RREADY),
    .m_axi_gmem_0_RDATA(m_axi_gmem_0_RDATA),
    .m_axi_gmem_0_RLAST(m_axi_gmem_0_RLAST),
    .m_axi_gmem_0_RID(m_axi_gmem_0_RID),
    .m_axi_gmem_0_RFIFONUM(m_axi_gmem_0_RFIFONUM),
    .m_axi_gmem_0_RUSER(m_axi_gmem_0_RUSER),
    .m_axi_gmem_0_RRESP(m_axi_gmem_0_RRESP),
    .m_axi_gmem_0_BVALID(1'b0),
    .m_axi_gmem_0_BREADY(grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_BREADY),
    .m_axi_gmem_0_BRESP(2'd0),
    .m_axi_gmem_0_BID(1'd0),
    .m_axi_gmem_0_BUSER(1'd0),
    .A_dram(A_dram_read_reg_311),
    .rows(rows_read_reg_306),
    .cols(cols_read_reg_301),
    .t_capacity(t_capacity_read_reg_296),
    .M_e_address0(grp_load_matrix_from_dram_safe_fu_174_M_e_address0),
    .M_e_ce0(grp_load_matrix_from_dram_safe_fu_174_M_e_ce0),
    .M_e_we0(grp_load_matrix_from_dram_safe_fu_174_M_e_we0),
    .M_e_d0(grp_load_matrix_from_dram_safe_fu_174_M_e_d0),
    .M_rows(grp_load_matrix_from_dram_safe_fu_174_M_rows),
    .M_rows_ap_vld(grp_load_matrix_from_dram_safe_fu_174_M_rows_ap_vld),
    .M_cols(grp_load_matrix_from_dram_safe_fu_174_M_cols),
    .M_cols_ap_vld(grp_load_matrix_from_dram_safe_fu_174_M_cols_ap_vld),
    .M_t(grp_load_matrix_from_dram_safe_fu_174_M_t),
    .M_t_ap_vld(grp_load_matrix_from_dram_safe_fu_174_M_t_ap_vld),
    .M_t_capacity(grp_load_matrix_from_dram_safe_fu_174_M_t_capacity),
    .M_t_capacity_ap_vld(grp_load_matrix_from_dram_safe_fu_174_M_t_capacity_ap_vld)
);

fmm_reduce_kernel_greedy_potential_reduce_with_debug grp_greedy_potential_reduce_with_debug_fu_198(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_greedy_potential_reduce_with_debug_fu_198_ap_start),
    .ap_done(grp_greedy_potential_reduce_with_debug_fu_198_ap_done),
    .ap_idle(grp_greedy_potential_reduce_with_debug_fu_198_ap_idle),
    .ap_ready(grp_greedy_potential_reduce_with_debug_fu_198_ap_ready),
    .k1(k1_read_reg_291),
    .k2(k2_read_reg_286),
    .m_axi_gmem2_0_AWVALID(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWVALID),
    .m_axi_gmem2_0_AWREADY(m_axi_gmem2_0_AWREADY),
    .m_axi_gmem2_0_AWADDR(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWADDR),
    .m_axi_gmem2_0_AWID(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWID),
    .m_axi_gmem2_0_AWLEN(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWLEN),
    .m_axi_gmem2_0_AWSIZE(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWSIZE),
    .m_axi_gmem2_0_AWBURST(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWBURST),
    .m_axi_gmem2_0_AWLOCK(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWLOCK),
    .m_axi_gmem2_0_AWCACHE(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWCACHE),
    .m_axi_gmem2_0_AWPROT(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWPROT),
    .m_axi_gmem2_0_AWQOS(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWQOS),
    .m_axi_gmem2_0_AWREGION(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWREGION),
    .m_axi_gmem2_0_AWUSER(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWUSER),
    .m_axi_gmem2_0_WVALID(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WVALID),
    .m_axi_gmem2_0_WREADY(m_axi_gmem2_0_WREADY),
    .m_axi_gmem2_0_WDATA(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WDATA),
    .m_axi_gmem2_0_WSTRB(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WSTRB),
    .m_axi_gmem2_0_WLAST(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WLAST),
    .m_axi_gmem2_0_WID(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WID),
    .m_axi_gmem2_0_WUSER(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WUSER),
    .m_axi_gmem2_0_ARVALID(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARVALID),
    .m_axi_gmem2_0_ARREADY(1'b0),
    .m_axi_gmem2_0_ARADDR(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARADDR),
    .m_axi_gmem2_0_ARID(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARID),
    .m_axi_gmem2_0_ARLEN(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARLEN),
    .m_axi_gmem2_0_ARSIZE(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARSIZE),
    .m_axi_gmem2_0_ARBURST(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARBURST),
    .m_axi_gmem2_0_ARLOCK(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARLOCK),
    .m_axi_gmem2_0_ARCACHE(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARCACHE),
    .m_axi_gmem2_0_ARPROT(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARPROT),
    .m_axi_gmem2_0_ARQOS(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARQOS),
    .m_axi_gmem2_0_ARREGION(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARREGION),
    .m_axi_gmem2_0_ARUSER(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_ARUSER),
    .m_axi_gmem2_0_RVALID(1'b0),
    .m_axi_gmem2_0_RREADY(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_RREADY),
    .m_axi_gmem2_0_RDATA(32'd0),
    .m_axi_gmem2_0_RLAST(1'b0),
    .m_axi_gmem2_0_RID(1'd0),
    .m_axi_gmem2_0_RFIFONUM(9'd0),
    .m_axi_gmem2_0_RUSER(1'd0),
    .m_axi_gmem2_0_RRESP(2'd0),
    .m_axi_gmem2_0_BVALID(m_axi_gmem2_0_BVALID),
    .m_axi_gmem2_0_BREADY(grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_BREADY),
    .m_axi_gmem2_0_BRESP(m_axi_gmem2_0_BRESP),
    .m_axi_gmem2_0_BID(m_axi_gmem2_0_BID),
    .m_axi_gmem2_0_BUSER(m_axi_gmem2_0_BUSER),
    .debug_dram(debug_dram_read_reg_280),
    .debug_capacity(debug_capacity_read_reg_275),
    .M_e_address0(grp_greedy_potential_reduce_with_debug_fu_198_M_e_address0),
    .M_e_ce0(grp_greedy_potential_reduce_with_debug_fu_198_M_e_ce0),
    .M_e_we0(grp_greedy_potential_reduce_with_debug_fu_198_M_e_we0),
    .M_e_d0(grp_greedy_potential_reduce_with_debug_fu_198_M_e_d0),
    .M_e_q0(M_e_q0),
    .M_e_address1(grp_greedy_potential_reduce_with_debug_fu_198_M_e_address1),
    .M_e_ce1(grp_greedy_potential_reduce_with_debug_fu_198_M_e_ce1),
    .M_e_we1(grp_greedy_potential_reduce_with_debug_fu_198_M_e_we1),
    .M_e_d1(grp_greedy_potential_reduce_with_debug_fu_198_M_e_d1),
    .M_e_q1(M_e_q1),
    .M_cols(M_cols),
    .M_rows(M_rows),
    .M_t_i(M_t),
    .M_t_o(grp_greedy_potential_reduce_with_debug_fu_198_M_t_o),
    .M_t_o_ap_vld(grp_greedy_potential_reduce_with_debug_fu_198_M_t_o_ap_vld),
    .M_t_capacity(M_t_capacity)
);

fmm_reduce_kernel_store_matrix_to_dram_safe grp_store_matrix_to_dram_safe_fu_218(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(grp_store_matrix_to_dram_safe_fu_218_ap_start),
    .ap_done(grp_store_matrix_to_dram_safe_fu_218_ap_done),
    .ap_idle(grp_store_matrix_to_dram_safe_fu_218_ap_idle),
    .ap_ready(grp_store_matrix_to_dram_safe_fu_218_ap_ready),
    .m_axi_gmem_0_AWVALID(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWVALID),
    .m_axi_gmem_0_AWREADY(m_axi_gmem_0_AWREADY),
    .m_axi_gmem_0_AWADDR(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWADDR),
    .m_axi_gmem_0_AWID(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWID),
    .m_axi_gmem_0_AWLEN(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWLEN),
    .m_axi_gmem_0_AWSIZE(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWSIZE),
    .m_axi_gmem_0_AWBURST(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWBURST),
    .m_axi_gmem_0_AWLOCK(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWLOCK),
    .m_axi_gmem_0_AWCACHE(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWCACHE),
    .m_axi_gmem_0_AWPROT(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWPROT),
    .m_axi_gmem_0_AWQOS(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWQOS),
    .m_axi_gmem_0_AWREGION(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWREGION),
    .m_axi_gmem_0_AWUSER(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWUSER),
    .m_axi_gmem_0_WVALID(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WVALID),
    .m_axi_gmem_0_WREADY(m_axi_gmem_0_WREADY),
    .m_axi_gmem_0_WDATA(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WDATA),
    .m_axi_gmem_0_WSTRB(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WSTRB),
    .m_axi_gmem_0_WLAST(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WLAST),
    .m_axi_gmem_0_WID(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WID),
    .m_axi_gmem_0_WUSER(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WUSER),
    .m_axi_gmem_0_ARVALID(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARVALID),
    .m_axi_gmem_0_ARREADY(1'b0),
    .m_axi_gmem_0_ARADDR(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARADDR),
    .m_axi_gmem_0_ARID(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARID),
    .m_axi_gmem_0_ARLEN(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARLEN),
    .m_axi_gmem_0_ARSIZE(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARSIZE),
    .m_axi_gmem_0_ARBURST(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARBURST),
    .m_axi_gmem_0_ARLOCK(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARLOCK),
    .m_axi_gmem_0_ARCACHE(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARCACHE),
    .m_axi_gmem_0_ARPROT(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARPROT),
    .m_axi_gmem_0_ARQOS(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARQOS),
    .m_axi_gmem_0_ARREGION(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARREGION),
    .m_axi_gmem_0_ARUSER(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_ARUSER),
    .m_axi_gmem_0_RVALID(1'b0),
    .m_axi_gmem_0_RREADY(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_RREADY),
    .m_axi_gmem_0_RDATA(32'd0),
    .m_axi_gmem_0_RLAST(1'b0),
    .m_axi_gmem_0_RID(1'd0),
    .m_axi_gmem_0_RFIFONUM(9'd0),
    .m_axi_gmem_0_RUSER(1'd0),
    .m_axi_gmem_0_RRESP(2'd0),
    .m_axi_gmem_0_BVALID(m_axi_gmem_0_BVALID),
    .m_axi_gmem_0_BREADY(grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_BREADY),
    .m_axi_gmem_0_BRESP(m_axi_gmem_0_BRESP),
    .m_axi_gmem_0_BID(m_axi_gmem_0_BID),
    .m_axi_gmem_0_BUSER(m_axi_gmem_0_BUSER),
    .A_dram(A_dram_read_reg_311),
    .M_rows(M_rows),
    .M_cols(M_cols),
    .M_e_address0(grp_store_matrix_to_dram_safe_fu_218_M_e_address0),
    .M_e_ce0(grp_store_matrix_to_dram_safe_fu_218_M_e_ce0),
    .M_e_q0(M_e_q0)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_state1;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_state8) & (1'b1 == ap_CS_fsm_state8))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_greedy_potential_reduce_with_debug_fu_198_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state10)) begin
            grp_greedy_potential_reduce_with_debug_fu_198_ap_start_reg <= 1'b1;
        end else if ((grp_greedy_potential_reduce_with_debug_fu_198_ap_ready == 1'b1)) begin
            grp_greedy_potential_reduce_with_debug_fu_198_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_load_matrix_from_dram_safe_fu_174_ap_start_reg <= 1'b0;
    end else begin
        if (((1'b0 == ap_block_state1_ignore_call0) & (1'd1 == and_ln307_fu_231_p2) & (1'b1 == ap_CS_fsm_state1))) begin
            grp_load_matrix_from_dram_safe_fu_174_ap_start_reg <= 1'b1;
        end else if ((grp_load_matrix_from_dram_safe_fu_174_ap_ready == 1'b1)) begin
            grp_load_matrix_from_dram_safe_fu_174_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        grp_store_matrix_to_dram_safe_fu_218_ap_start_reg <= 1'b0;
    end else begin
        if ((1'b1 == ap_CS_fsm_state12)) begin
            grp_store_matrix_to_dram_safe_fu_218_ap_start_reg <= 1'b1;
        end else if ((grp_store_matrix_to_dram_safe_fu_218_ap_ready == 1'b1)) begin
            grp_store_matrix_to_dram_safe_fu_218_ap_start_reg <= 1'b0;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((grp_greedy_potential_reduce_with_debug_fu_198_M_t_o_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state11))) begin
        M_t <= grp_greedy_potential_reduce_with_debug_fu_198_M_t_o;
    end else if (((grp_load_matrix_from_dram_safe_fu_174_M_t_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state9))) begin
        M_t <= grp_load_matrix_from_dram_safe_fu_174_M_t;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1))) begin
        A_dram_read_reg_311 <= A_dram_dout;
        and_ln307_reg_317 <= and_ln307_fu_231_p2;
        cols_read_reg_301 <= cols_dout;
        debug_capacity_read_reg_275 <= debug_capacity_dout;
        debug_dram_read_reg_280 <= debug_dram_dout;
        icmp_ln308_reg_321 <= icmp_ln308_fu_237_p2;
        k1_read_reg_291 <= k1_dout;
        k2_read_reg_286 <= k2_dout;
        p_read_2_reg_270 <= p_read;
        rows_read_reg_306 <= rows_dout;
        t_capacity_read_reg_296 <= t_capacity_dout;
    end
end

always @ (posedge ap_clk) begin
    if (((grp_load_matrix_from_dram_safe_fu_174_M_cols_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state9))) begin
        M_cols <= grp_load_matrix_from_dram_safe_fu_174_M_cols;
    end
end

always @ (posedge ap_clk) begin
    if (((grp_load_matrix_from_dram_safe_fu_174_M_rows_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state9))) begin
        M_rows <= grp_load_matrix_from_dram_safe_fu_174_M_rows;
    end
end

always @ (posedge ap_clk) begin
    if (((grp_load_matrix_from_dram_safe_fu_174_M_t_capacity_ap_vld == 1'b1) & (1'b1 == ap_CS_fsm_state9))) begin
        M_t_capacity <= grp_load_matrix_from_dram_safe_fu_174_M_t_capacity;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_state2) & (m_axi_gmem2_0_AWREADY == 1'b1))) begin
        select_ln309_reg_325[2 : 0] <= select_ln309_fu_243_p3[2 : 0];
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        A_dram_blk_n = A_dram_empty_n;
    end else begin
        A_dram_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1))) begin
        A_dram_read = 1'b1;
    end else begin
        A_dram_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        M_e_address0 = grp_store_matrix_to_dram_safe_fu_218_M_e_address0;
    end else if ((1'b1 == ap_CS_fsm_state11)) begin
        M_e_address0 = grp_greedy_potential_reduce_with_debug_fu_198_M_e_address0;
    end else if ((1'b1 == ap_CS_fsm_state9)) begin
        M_e_address0 = grp_load_matrix_from_dram_safe_fu_174_M_e_address0;
    end else begin
        M_e_address0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state13)) begin
        M_e_ce0 = grp_store_matrix_to_dram_safe_fu_218_M_e_ce0;
    end else if ((1'b1 == ap_CS_fsm_state11)) begin
        M_e_ce0 = grp_greedy_potential_reduce_with_debug_fu_198_M_e_ce0;
    end else if ((1'b1 == ap_CS_fsm_state9)) begin
        M_e_ce0 = grp_load_matrix_from_dram_safe_fu_174_M_e_ce0;
    end else begin
        M_e_ce0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state11)) begin
        M_e_ce1 = grp_greedy_potential_reduce_with_debug_fu_198_M_e_ce1;
    end else begin
        M_e_ce1 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state11)) begin
        M_e_d0 = grp_greedy_potential_reduce_with_debug_fu_198_M_e_d0;
    end else if ((1'b1 == ap_CS_fsm_state9)) begin
        M_e_d0 = grp_load_matrix_from_dram_safe_fu_174_M_e_d0;
    end else begin
        M_e_d0 = 'bx;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state11)) begin
        M_e_we0 = grp_greedy_potential_reduce_with_debug_fu_198_M_e_we0;
    end else if ((1'b1 == ap_CS_fsm_state9)) begin
        M_e_we0 = grp_load_matrix_from_dram_safe_fu_174_M_e_we0;
    end else begin
        M_e_we0 = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state11)) begin
        M_e_we1 = grp_greedy_potential_reduce_with_debug_fu_198_M_e_we1;
    end else begin
        M_e_we1 = 1'b0;
    end
end

assign ap_ST_fsm_state10_blk = 1'b0;

always @ (*) begin
    if ((grp_greedy_potential_reduce_with_debug_fu_198_ap_done == 1'b0)) begin
        ap_ST_fsm_state11_blk = 1'b1;
    end else begin
        ap_ST_fsm_state11_blk = 1'b0;
    end
end

assign ap_ST_fsm_state12_blk = 1'b0;

always @ (*) begin
    if ((grp_store_matrix_to_dram_safe_fu_218_ap_done == 1'b0)) begin
        ap_ST_fsm_state13_blk = 1'b1;
    end else begin
        ap_ST_fsm_state13_blk = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_block_state1)) begin
        ap_ST_fsm_state1_blk = 1'b1;
    end else begin
        ap_ST_fsm_state1_blk = 1'b0;
    end
end

always @ (*) begin
    if ((m_axi_gmem2_0_AWREADY == 1'b0)) begin
        ap_ST_fsm_state2_blk = 1'b1;
    end else begin
        ap_ST_fsm_state2_blk = 1'b0;
    end
end

always @ (*) begin
    if ((m_axi_gmem2_0_WREADY == 1'b0)) begin
        ap_ST_fsm_state3_blk = 1'b1;
    end else begin
        ap_ST_fsm_state3_blk = 1'b0;
    end
end

assign ap_ST_fsm_state4_blk = 1'b0;

assign ap_ST_fsm_state5_blk = 1'b0;

assign ap_ST_fsm_state6_blk = 1'b0;

assign ap_ST_fsm_state7_blk = 1'b0;

always @ (*) begin
    if ((1'b1 == ap_block_state8)) begin
        ap_ST_fsm_state8_blk = 1'b1;
    end else begin
        ap_ST_fsm_state8_blk = 1'b0;
    end
end

always @ (*) begin
    if ((grp_load_matrix_from_dram_safe_fu_174_ap_done == 1'b0)) begin
        ap_ST_fsm_state9_blk = 1'b1;
    end else begin
        ap_ST_fsm_state9_blk = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state8) & (1'b1 == ap_CS_fsm_state8))) begin
        ap_done = 1'b1;
    end else begin
        ap_done = ap_done_reg;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state1) & (ap_start == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state8) & (1'b1 == ap_CS_fsm_state8))) begin
        ap_ready = 1'b1;
    end else begin
        ap_ready = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        cols_blk_n = cols_empty_n;
    end else begin
        cols_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1))) begin
        cols_read = 1'b1;
    end else begin
        cols_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        debug_capacity_blk_n = debug_capacity_empty_n;
    end else begin
        debug_capacity_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1))) begin
        debug_capacity_read = 1'b1;
    end else begin
        debug_capacity_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        debug_dram_blk_n = debug_dram_empty_n;
    end else begin
        debug_dram_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1))) begin
        debug_dram_read = 1'b1;
    end else begin
        debug_dram_read = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state2)) begin
        gmem2_blk_n_AW = m_axi_gmem2_0_AWREADY;
    end else begin
        gmem2_blk_n_AW = 1'b1;
    end
end

always @ (*) begin
    if (((icmp_ln308_reg_321 == 1'd1) & (1'b1 == ap_CS_fsm_state8) & (1'd0 == and_ln307_reg_317))) begin
        gmem2_blk_n_B = m_axi_gmem2_0_BVALID;
    end else begin
        gmem2_blk_n_B = 1'b1;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        gmem2_blk_n_W = m_axi_gmem2_0_WREADY;
    end else begin
        gmem2_blk_n_W = 1'b1;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        k1_blk_n = k1_empty_n;
    end else begin
        k1_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1))) begin
        k1_read = 1'b1;
    end else begin
        k1_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        k2_blk_n = k2_empty_n;
    end else begin
        k2_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1))) begin
        k2_read = 1'b1;
    end else begin
        k2_read = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) & (m_axi_gmem2_0_AWREADY == 1'b1))) begin
        m_axi_gmem2_0_AWADDR = sext_ln309_fu_259_p1;
    end else if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWADDR = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWADDR;
    end else begin
        m_axi_gmem2_0_AWADDR = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWBURST = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWBURST;
    end else begin
        m_axi_gmem2_0_AWBURST = 2'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWCACHE = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWCACHE;
    end else begin
        m_axi_gmem2_0_AWCACHE = 4'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWID = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWID;
    end else begin
        m_axi_gmem2_0_AWID = 1'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) & (m_axi_gmem2_0_AWREADY == 1'b1))) begin
        m_axi_gmem2_0_AWLEN = 64'd1;
    end else if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWLEN = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWLEN;
    end else begin
        m_axi_gmem2_0_AWLEN = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWLOCK = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWLOCK;
    end else begin
        m_axi_gmem2_0_AWLOCK = 2'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWPROT = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWPROT;
    end else begin
        m_axi_gmem2_0_AWPROT = 3'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWQOS = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWQOS;
    end else begin
        m_axi_gmem2_0_AWQOS = 4'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWREGION = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWREGION;
    end else begin
        m_axi_gmem2_0_AWREGION = 4'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWSIZE = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWSIZE;
    end else begin
        m_axi_gmem2_0_AWSIZE = 3'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWUSER = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWUSER;
    end else begin
        m_axi_gmem2_0_AWUSER = 1'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state2) & (m_axi_gmem2_0_AWREADY == 1'b1))) begin
        m_axi_gmem2_0_AWVALID = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_AWVALID = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_AWVALID;
    end else begin
        m_axi_gmem2_0_AWVALID = 1'b0;
    end
end

always @ (*) begin
    if (((ap_predicate_op49_writeresp_state8 == 1'b1) & (1'b0 == ap_block_state8) & (1'b1 == ap_CS_fsm_state8))) begin
        m_axi_gmem2_0_BREADY = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_BREADY = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_BREADY;
    end else begin
        m_axi_gmem2_0_BREADY = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        m_axi_gmem2_0_WDATA = select_ln309_reg_325;
    end else if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_WDATA = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WDATA;
    end else begin
        m_axi_gmem2_0_WDATA = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_WID = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WID;
    end else begin
        m_axi_gmem2_0_WID = 1'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_WLAST = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WLAST;
    end else begin
        m_axi_gmem2_0_WLAST = 1'b0;
    end
end

always @ (*) begin
    if ((1'b1 == ap_CS_fsm_state3)) begin
        m_axi_gmem2_0_WSTRB = 4'd15;
    end else if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_WSTRB = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WSTRB;
    end else begin
        m_axi_gmem2_0_WSTRB = 'bx;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_WUSER = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WUSER;
    end else begin
        m_axi_gmem2_0_WUSER = 1'd0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state3) & (m_axi_gmem2_0_WREADY == 1'b1))) begin
        m_axi_gmem2_0_WVALID = 1'b1;
    end else if (((1'b1 == ap_CS_fsm_state11) | (1'b1 == ap_CS_fsm_state10))) begin
        m_axi_gmem2_0_WVALID = grp_greedy_potential_reduce_with_debug_fu_198_m_axi_gmem2_0_WVALID;
    end else begin
        m_axi_gmem2_0_WVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state1))) begin
        m_axi_gmem_0_ARVALID = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARVALID;
    end else begin
        m_axi_gmem_0_ARVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        m_axi_gmem_0_AWVALID = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWVALID;
    end else begin
        m_axi_gmem_0_AWVALID = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        m_axi_gmem_0_BREADY = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_BREADY;
    end else begin
        m_axi_gmem_0_BREADY = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state9) | (1'b1 == ap_CS_fsm_state1))) begin
        m_axi_gmem_0_RREADY = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_RREADY;
    end else begin
        m_axi_gmem_0_RREADY = 1'b0;
    end
end

always @ (*) begin
    if (((1'b1 == ap_CS_fsm_state13) | (1'b1 == ap_CS_fsm_state12))) begin
        m_axi_gmem_0_WVALID = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WVALID;
    end else begin
        m_axi_gmem_0_WVALID = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        rows_blk_n = rows_empty_n;
    end else begin
        rows_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1))) begin
        rows_read = 1'b1;
    end else begin
        rows_read = 1'b0;
    end
end

always @ (*) begin
    if ((~((ap_done_reg == 1'b1) | (ap_start == 1'b0)) & (1'b1 == ap_CS_fsm_state1))) begin
        t_capacity_blk_n = t_capacity_empty_n;
    end else begin
        t_capacity_blk_n = 1'b1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1))) begin
        t_capacity_read = 1'b1;
    end else begin
        t_capacity_read = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_state1 : begin
            if (((icmp_ln308_fu_237_p2 == 1'd0) & (1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1) & (1'd0 == and_ln307_fu_231_p2))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else if (((icmp_ln308_fu_237_p2 == 1'd1) & (1'b0 == ap_block_state1) & (1'b1 == ap_CS_fsm_state1) & (1'd0 == and_ln307_fu_231_p2))) begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end else if (((1'b0 == ap_block_state1) & (1'd1 == and_ln307_fu_231_p2) & (1'b1 == ap_CS_fsm_state1))) begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end
        end
        ap_ST_fsm_state2 : begin
            if (((1'b1 == ap_CS_fsm_state2) & (m_axi_gmem2_0_AWREADY == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state2;
            end
        end
        ap_ST_fsm_state3 : begin
            if (((1'b1 == ap_CS_fsm_state3) & (m_axi_gmem2_0_WREADY == 1'b1))) begin
                ap_NS_fsm = ap_ST_fsm_state4;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state3;
            end
        end
        ap_ST_fsm_state4 : begin
            ap_NS_fsm = ap_ST_fsm_state5;
        end
        ap_ST_fsm_state5 : begin
            ap_NS_fsm = ap_ST_fsm_state6;
        end
        ap_ST_fsm_state6 : begin
            ap_NS_fsm = ap_ST_fsm_state7;
        end
        ap_ST_fsm_state7 : begin
            ap_NS_fsm = ap_ST_fsm_state8;
        end
        ap_ST_fsm_state8 : begin
            if (((1'b0 == ap_block_state8) & (1'b1 == ap_CS_fsm_state8))) begin
                ap_NS_fsm = ap_ST_fsm_state1;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end
        end
        ap_ST_fsm_state9 : begin
            if (((grp_load_matrix_from_dram_safe_fu_174_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state9))) begin
                ap_NS_fsm = ap_ST_fsm_state10;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state9;
            end
        end
        ap_ST_fsm_state10 : begin
            ap_NS_fsm = ap_ST_fsm_state11;
        end
        ap_ST_fsm_state11 : begin
            if (((grp_greedy_potential_reduce_with_debug_fu_198_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state11))) begin
                ap_NS_fsm = ap_ST_fsm_state12;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state11;
            end
        end
        ap_ST_fsm_state12 : begin
            ap_NS_fsm = ap_ST_fsm_state13;
        end
        ap_ST_fsm_state13 : begin
            if (((grp_store_matrix_to_dram_safe_fu_218_ap_done == 1'b1) & (1'b1 == ap_CS_fsm_state13))) begin
                ap_NS_fsm = ap_ST_fsm_state8;
            end else begin
                ap_NS_fsm = ap_ST_fsm_state13;
            end
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign and_ln307_fu_231_p2 = (p_read1 & p_read);

assign ap_CS_fsm_state1 = ap_CS_fsm[32'd0];

assign ap_CS_fsm_state10 = ap_CS_fsm[32'd9];

assign ap_CS_fsm_state11 = ap_CS_fsm[32'd10];

assign ap_CS_fsm_state12 = ap_CS_fsm[32'd11];

assign ap_CS_fsm_state13 = ap_CS_fsm[32'd12];

assign ap_CS_fsm_state2 = ap_CS_fsm[32'd1];

assign ap_CS_fsm_state3 = ap_CS_fsm[32'd2];

assign ap_CS_fsm_state8 = ap_CS_fsm[32'd7];

assign ap_CS_fsm_state9 = ap_CS_fsm[32'd8];

always @ (*) begin
    ap_block_state1 = ((rows_empty_n == 1'b0) | (1'b0 == A_dram_empty_n) | (ap_done_reg == 1'b1) | (debug_capacity_empty_n == 1'b0) | (ap_start == 1'b0) | (debug_dram_empty_n == 1'b0) | (k2_empty_n == 1'b0) | (k1_empty_n == 1'b0) | (t_capacity_empty_n == 1'b0) | (cols_empty_n == 1'b0));
end

always @ (*) begin
    ap_block_state1_ignore_call0 = ((rows_empty_n == 1'b0) | (1'b0 == A_dram_empty_n) | (ap_done_reg == 1'b1) | (debug_capacity_empty_n == 1'b0) | (ap_start == 1'b0) | (debug_dram_empty_n == 1'b0) | (k2_empty_n == 1'b0) | (k1_empty_n == 1'b0) | (t_capacity_empty_n == 1'b0) | (cols_empty_n == 1'b0));
end

always @ (*) begin
    ap_block_state8 = ((ap_predicate_op49_writeresp_state8 == 1'b1) & (m_axi_gmem2_0_BVALID == 1'b0));
end

always @ (*) begin
    ap_predicate_op49_writeresp_state8 = ((icmp_ln308_reg_321 == 1'd1) & (1'd0 == and_ln307_reg_317));
end

assign grp_greedy_potential_reduce_with_debug_fu_198_ap_start = grp_greedy_potential_reduce_with_debug_fu_198_ap_start_reg;

assign grp_load_matrix_from_dram_safe_fu_174_ap_start = grp_load_matrix_from_dram_safe_fu_174_ap_start_reg;

assign grp_store_matrix_to_dram_safe_fu_218_ap_start = grp_store_matrix_to_dram_safe_fu_218_ap_start_reg;

assign icmp_ln308_fu_237_p2 = (($signed(debug_capacity_dout) > $signed(32'd0)) ? 1'b1 : 1'b0);

assign m_axi_gmem2_0_ARADDR = 64'd0;

assign m_axi_gmem2_0_ARBURST = 2'd0;

assign m_axi_gmem2_0_ARCACHE = 4'd0;

assign m_axi_gmem2_0_ARID = 1'd0;

assign m_axi_gmem2_0_ARLEN = 32'd0;

assign m_axi_gmem2_0_ARLOCK = 2'd0;

assign m_axi_gmem2_0_ARPROT = 3'd0;

assign m_axi_gmem2_0_ARQOS = 4'd0;

assign m_axi_gmem2_0_ARREGION = 4'd0;

assign m_axi_gmem2_0_ARSIZE = 3'd0;

assign m_axi_gmem2_0_ARUSER = 1'd0;

assign m_axi_gmem2_0_ARVALID = 1'b0;

assign m_axi_gmem2_0_RREADY = 1'b0;

assign m_axi_gmem_0_ARADDR = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARADDR;

assign m_axi_gmem_0_ARBURST = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARBURST;

assign m_axi_gmem_0_ARCACHE = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARCACHE;

assign m_axi_gmem_0_ARID = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARID;

assign m_axi_gmem_0_ARLEN = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARLEN;

assign m_axi_gmem_0_ARLOCK = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARLOCK;

assign m_axi_gmem_0_ARPROT = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARPROT;

assign m_axi_gmem_0_ARQOS = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARQOS;

assign m_axi_gmem_0_ARREGION = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARREGION;

assign m_axi_gmem_0_ARSIZE = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARSIZE;

assign m_axi_gmem_0_ARUSER = grp_load_matrix_from_dram_safe_fu_174_m_axi_gmem_0_ARUSER;

assign m_axi_gmem_0_AWADDR = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWADDR;

assign m_axi_gmem_0_AWBURST = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWBURST;

assign m_axi_gmem_0_AWCACHE = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWCACHE;

assign m_axi_gmem_0_AWID = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWID;

assign m_axi_gmem_0_AWLEN = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWLEN;

assign m_axi_gmem_0_AWLOCK = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWLOCK;

assign m_axi_gmem_0_AWPROT = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWPROT;

assign m_axi_gmem_0_AWQOS = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWQOS;

assign m_axi_gmem_0_AWREGION = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWREGION;

assign m_axi_gmem_0_AWSIZE = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWSIZE;

assign m_axi_gmem_0_AWUSER = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_AWUSER;

assign m_axi_gmem_0_WDATA = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WDATA;

assign m_axi_gmem_0_WID = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WID;

assign m_axi_gmem_0_WLAST = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WLAST;

assign m_axi_gmem_0_WSTRB = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WSTRB;

assign m_axi_gmem_0_WUSER = grp_store_matrix_to_dram_safe_fu_218_m_axi_gmem_0_WUSER;

assign select_ln309_fu_243_p3 = ((p_read_2_reg_270[0:0] == 1'b1) ? 32'd4294966395 : 32'd4294966396);

assign sext_ln309_fu_259_p1 = $signed(trunc_ln_fu_250_p4);

assign trunc_ln_fu_250_p4 = {{debug_dram_read_reg_280[63:2]}};

always @ (posedge ap_clk) begin
    select_ln309_reg_325[31:3] <= 29'b11111111111111111111110001111;
end

endmodule //fmm_reduce_kernel_Block_entry_proc
