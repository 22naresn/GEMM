`timescale 1 ns / 1 ps 

module fmm_reduce_kernel_greedy_potential_reduce_with_debug_Pipeline_VITIS_LOOP_163_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        zext_ln163,
        idxprom4_i12_i332_i_i,
        M_e_address0,
        M_e_ce0,
        M_e_q0,
        sext_ln163,
        move_type_1_out,
        move_type_1_out_ap_vld,
        row2_1_out,
        row2_1_out_ap_vld
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [31:0] zext_ln163;
input  [16:0] idxprom4_i12_i332_i_i;
output  [16:0] M_e_address0;
output   M_e_ce0;
input  [31:0] M_e_q0;
input  [31:0] sext_ln163;
output  [31:0] move_type_1_out;
output   move_type_1_out_ap_vld;
output  [31:0] row2_1_out;
output   row2_1_out_ap_vld;

reg ap_idle;
reg move_type_1_out_ap_vld;
reg row2_1_out_ap_vld;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_idle_pp0;
wire    ap_block_pp0_stage0_subdone;
wire   [0:0] or_cond284_i_fu_219_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire    ap_block_pp0_stage0_11001;
wire   [31:0] trunc_ln166_fu_174_p1;
reg   [31:0] trunc_ln166_reg_264;
wire   [33:0] add_ln163_fu_178_p2;
reg   [33:0] add_ln163_reg_269;
wire   [0:0] icmp_ln163_fu_184_p2;
reg   [0:0] icmp_ln163_reg_274;
wire   [63:0] zext_ln165_fu_169_p1;
wire    ap_block_pp0_stage0;
reg   [31:0] move_type_fu_46;
wire   [31:0] move_type_4_fu_202_p3;
wire    ap_loop_init;
reg   [31:0] row2_fu_50;
wire   [31:0] row2_4_fu_211_p3;
reg   [33:0] r_fu_54;
wire   [33:0] zext_ln163_cast_fu_107_p1;
reg   [33:0] ap_sig_allocacmp_r_2;
wire    ap_block_pp0_stage0_01001;
reg    M_e_ce0_local;
wire   [26:0] trunc_ln165_fu_129_p1;
wire   [28:0] trunc_ln165_3_fu_141_p1;
wire   [34:0] p_shl_fu_133_p3;
wire   [34:0] p_shl6_fu_145_p3;
wire   [34:0] add_ln165_2_fu_153_p2;
wire   [16:0] trunc_ln165_4_fu_159_p1;
wire   [16:0] add_ln165_fu_163_p2;
wire  signed [33:0] sext_ln163_cast_fu_103_p1;
wire   [0:0] icmp_ln166_fu_196_p2;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ready_sig;
wire    ap_done_sig;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 move_type_fu_46 = 32'd0;
#0 row2_fu_50 = 32'd0;
#0 r_fu_54 = 34'd0;
#0 ap_done_reg = 1'b0;
end

fmm_reduce_kernel_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready_sig),
    .ap_done(ap_done_sig),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            move_type_fu_46 <= 32'd0;
        end else if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            move_type_fu_46 <= move_type_4_fu_202_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            r_fu_54 <= zext_ln163_cast_fu_107_p1;
        end else if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            r_fu_54 <= add_ln163_reg_269;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            row2_fu_50 <= 32'd4294967295;
        end else if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            row2_fu_50 <= row2_4_fu_211_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln163_reg_269 <= add_ln163_fu_178_p2;
        icmp_ln163_reg_274 <= icmp_ln163_fu_184_p2;
        trunc_ln166_reg_264 <= trunc_ln166_fu_174_p1;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        M_e_ce0_local = 1'b1;
    end else begin
        M_e_ce0_local = 1'b0;
    end
end

always @ (*) begin
    if (((or_cond284_i_fu_219_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            ap_sig_allocacmp_r_2 = zext_ln163_cast_fu_107_p1;
        end else if ((ap_enable_reg_pp0_iter1 == 1'b1)) begin
            ap_sig_allocacmp_r_2 = add_ln163_reg_269;
        end else begin
            ap_sig_allocacmp_r_2 = r_fu_54;
        end
    end else begin
        ap_sig_allocacmp_r_2 = r_fu_54;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready == 1'b1) & (or_cond284_i_fu_219_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        move_type_1_out_ap_vld = 1'b1;
    end else begin
        move_type_1_out_ap_vld = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready == 1'b1) & (or_cond284_i_fu_219_p2 == 1'd0) & (1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        row2_1_out_ap_vld = 1'b1;
    end else begin
        row2_1_out_ap_vld = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign M_e_address0 = zext_ln165_fu_169_p1;

assign M_e_ce0 = M_e_ce0_local;

assign add_ln163_fu_178_p2 = ($signed(ap_sig_allocacmp_r_2) + $signed(34'd17179869183));

assign add_ln165_2_fu_153_p2 = (p_shl_fu_133_p3 + p_shl6_fu_145_p3);

assign add_ln165_fu_163_p2 = (trunc_ln165_4_fu_159_p1 + idxprom4_i12_i332_i_i);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_done = ap_done_sig;

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign ap_ready = ap_ready_sig;

assign icmp_ln163_fu_184_p2 = (($signed(add_ln163_fu_178_p2) > $signed(sext_ln163_cast_fu_103_p1)) ? 1'b1 : 1'b0);

assign icmp_ln166_fu_196_p2 = ((M_e_q0 == 32'd0) ? 1'b1 : 1'b0);

assign move_type_1_out = ((icmp_ln166_fu_196_p2[0:0] == 1'b1) ? move_type_fu_46 : M_e_q0);

assign move_type_4_fu_202_p3 = ((icmp_ln166_fu_196_p2[0:0] == 1'b1) ? move_type_fu_46 : M_e_q0);

assign or_cond284_i_fu_219_p2 = (icmp_ln166_fu_196_p2 & icmp_ln163_reg_274);

assign p_shl6_fu_145_p3 = {{trunc_ln165_3_fu_141_p1}, {6'd0}};

assign p_shl_fu_133_p3 = {{trunc_ln165_fu_129_p1}, {8'd0}};

assign row2_1_out = ((icmp_ln166_fu_196_p2[0:0] == 1'b1) ? row2_fu_50 : trunc_ln166_reg_264);

assign row2_4_fu_211_p3 = ((icmp_ln166_fu_196_p2[0:0] == 1'b1) ? row2_fu_50 : trunc_ln166_reg_264);

assign sext_ln163_cast_fu_103_p1 = $signed(sext_ln163);

assign trunc_ln165_3_fu_141_p1 = ap_sig_allocacmp_r_2[28:0];

assign trunc_ln165_4_fu_159_p1 = add_ln165_2_fu_153_p2[16:0];

assign trunc_ln165_fu_129_p1 = ap_sig_allocacmp_r_2[26:0];

assign trunc_ln166_fu_174_p1 = ap_sig_allocacmp_r_2[31:0];

assign zext_ln163_cast_fu_107_p1 = zext_ln163;

assign zext_ln165_fu_169_p1 = add_ln165_fu_163_p2;

endmodule //fmm_reduce_kernel_greedy_potential_reduce_with_debug_Pipeline_VITIS_LOOP_163_2
