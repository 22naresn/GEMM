`timescale 1 ns / 1 ps 

module fmm_reduce_kernel_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        M_e_address0,
        M_e_ce0,
        M_e_we0,
        M_e_d0
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output  [16:0] M_e_address0;
output   M_e_ce0;
output   M_e_we0;
output  [31:0] M_e_d0;

reg ap_idle;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_idle_pp0;
wire    ap_block_pp0_stage0_subdone;
wire   [0:0] icmp_ln49_fu_84_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire   [16:0] add_ln53_fu_160_p2;
reg   [16:0] add_ln53_reg_215;
wire    ap_block_pp0_stage0_11001;
wire   [63:0] zext_ln53_1_fu_187_p1;
wire    ap_block_pp0_stage0;
reg   [8:0] c_fu_40;
wire   [8:0] add_ln51_fu_166_p2;
wire    ap_loop_init;
reg   [8:0] r_fu_44;
wire   [8:0] select_ln49_1_fu_122_p3;
reg   [16:0] indvar_flatten_fu_48;
wire   [16:0] add_ln49_1_fu_90_p2;
reg    M_e_we0_local;
reg    M_e_ce0_local;
wire   [0:0] icmp_ln51_fu_108_p2;
wire   [8:0] add_ln49_fu_102_p2;
wire   [14:0] tmp_1_fu_138_p3;
wire   [16:0] tmp_fu_130_p3;
wire   [16:0] zext_ln51_fu_146_p1;
wire   [8:0] select_ln49_fu_114_p3;
wire   [16:0] add_ln51_1_fu_150_p2;
wire   [16:0] zext_ln53_fu_156_p1;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ready_sig;
wire    ap_done_sig;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 c_fu_40 = 9'd0;
#0 r_fu_44 = 9'd0;
#0 indvar_flatten_fu_48 = 17'd0;
#0 ap_done_reg = 1'b0;
end

fmm_reduce_kernel_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready_sig),
    .ap_done(ap_done_sig),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            c_fu_40 <= 9'd0;
        end else if (((icmp_ln49_fu_84_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            c_fu_40 <= add_ln51_fu_166_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            indvar_flatten_fu_48 <= 17'd0;
        end else if (((icmp_ln49_fu_84_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            indvar_flatten_fu_48 <= add_ln49_1_fu_90_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            r_fu_44 <= 9'd0;
        end else if (((icmp_ln49_fu_84_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            r_fu_44 <= select_ln49_1_fu_122_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        add_ln53_reg_215 <= add_ln53_fu_160_p2;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        M_e_ce0_local = 1'b1;
    end else begin
        M_e_ce0_local = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        M_e_we0_local = 1'b1;
    end else begin
        M_e_we0_local = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln49_fu_84_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (ap_start_int == 1'b0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign M_e_address0 = zext_ln53_1_fu_187_p1;

assign M_e_ce0 = M_e_ce0_local;

assign M_e_d0 = 32'd0;

assign M_e_we0 = M_e_we0_local;

assign add_ln49_1_fu_90_p2 = (indvar_flatten_fu_48 + 17'd1);

assign add_ln49_fu_102_p2 = (r_fu_44 + 9'd1);

assign add_ln51_1_fu_150_p2 = (tmp_fu_130_p3 + zext_ln51_fu_146_p1);

assign add_ln51_fu_166_p2 = (select_ln49_fu_114_p3 + 9'd1);

assign add_ln53_fu_160_p2 = (add_ln51_1_fu_150_p2 + zext_ln53_fu_156_p1);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_done = ap_done_sig;

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign ap_ready = ap_ready_sig;

assign icmp_ln49_fu_84_p2 = ((indvar_flatten_fu_48 == 17'd102400) ? 1'b1 : 1'b0);

assign icmp_ln51_fu_108_p2 = ((c_fu_40 == 9'd320) ? 1'b1 : 1'b0);

assign select_ln49_1_fu_122_p3 = ((icmp_ln51_fu_108_p2[0:0] == 1'b1) ? add_ln49_fu_102_p2 : r_fu_44);

assign select_ln49_fu_114_p3 = ((icmp_ln51_fu_108_p2[0:0] == 1'b1) ? 9'd0 : c_fu_40);

assign tmp_1_fu_138_p3 = {{select_ln49_1_fu_122_p3}, {6'd0}};

assign tmp_fu_130_p3 = {{select_ln49_1_fu_122_p3}, {8'd0}};

assign zext_ln51_fu_146_p1 = tmp_1_fu_138_p3;

assign zext_ln53_1_fu_187_p1 = add_ln53_reg_215;

assign zext_ln53_fu_156_p1 = select_ln49_fu_114_p3;

endmodule //fmm_reduce_kernel_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_49_1_VITIS_LOOP_51_2
