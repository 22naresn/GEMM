`timescale 1 ns / 1 ps 

module fmm_reduce_kernel_greedy_potential_reduce_with_debug_Pipeline_VITIS_LOOP_192_2_VITIS_LOOP_115_1 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        zext_ln192,
        s_4,
        cols_non_t,
        mul_ln191,
        mul_ln117_1,
        M_e_address0,
        M_e_ce0,
        M_e_q0,
        M_e_address1,
        M_e_ce1,
        M_e_q1,
        s_9_out,
        s_9_out_ap_vld
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
input  [30:0] zext_ln192;
input  [31:0] s_4;
input  [31:0] cols_non_t;
input  [94:0] mul_ln191;
input  [16:0] mul_ln117_1;
output  [16:0] M_e_address0;
output   M_e_ce0;
input  [31:0] M_e_q0;
output  [16:0] M_e_address1;
output   M_e_ce1;
input  [31:0] M_e_q1;
output  [31:0] s_9_out;
output   s_9_out_ap_vld;

reg ap_idle;
reg s_9_out_ap_vld;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_idle_pp0;
wire    ap_block_pp0_stage0_subdone;
wire   [0:0] icmp_ln192_fu_201_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
wire    ap_block_pp0_stage0_11001;
wire   [0:0] icmp_ln115_fu_196_p2;
reg   [0:0] icmp_ln115_reg_582;
reg   [0:0] icmp_ln115_reg_582_pp0_iter2_reg;
reg   [0:0] icmp_ln192_reg_589;
reg   [0:0] icmp_ln192_reg_589_pp0_iter2_reg;
wire   [8:0] trunc_ln119_fu_237_p1;
reg   [8:0] trunc_ln119_reg_593;
wire   [10:0] trunc_ln119_2_fu_241_p1;
reg   [10:0] trunc_ln119_2_reg_598;
wire   [16:0] trunc_ln117_fu_245_p1;
reg   [16:0] trunc_ln117_reg_603;
wire   [63:0] zext_ln117_fu_294_p1;
wire    ap_block_pp0_stage0;
wire   [63:0] zext_ln119_fu_304_p1;
reg   [31:0] n_3_fu_66;
wire   [31:0] n_5_fu_482_p3;
wire    ap_loop_init;
reg   [31:0] p_fu_70;
wire   [31:0] p_6_fu_502_p3;
reg   [30:0] c_fu_74;
wire   [30:0] add_ln115_fu_249_p2;
reg   [31:0] s_5_fu_78;
wire   [31:0] select_ln192_1_fu_405_p3;
reg   [63:0] j_fu_82;
wire   [63:0] select_ln192_fu_229_p3;
wire   [63:0] zext_ln192_cast_fu_152_p1;
reg   [94:0] indvar_flatten8_fu_86;
wire   [94:0] add_ln192_fu_206_p2;
wire   [31:0] s_9_fu_382_p3;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
wire    ap_block_pp0_stage0_01001;
reg    M_e_ce1_local;
reg    M_e_ce0_local;
wire   [31:0] zext_ln115_fu_192_p1;
wire   [63:0] add_ln192_1_fu_215_p2;
wire   [30:0] select_ln193_fu_221_p3;
wire   [16:0] p_shl_fu_270_p3;
wire   [16:0] p_shl4_fu_277_p3;
wire   [16:0] add_ln117_fu_290_p2;
wire   [16:0] add_ln119_fu_284_p2;
wire   [16:0] add_ln119_2_fu_299_p2;
wire   [30:0] tmp_fu_318_p4;
wire   [31:0] add_ln196_fu_334_p2;
wire   [0:0] icmp_ln196_fu_328_p2;
wire   [31:0] s_6_fu_340_p2;
wire   [30:0] tmp_3_fu_354_p4;
wire   [31:0] s_7_fu_346_p3;
wire   [31:0] add_ln197_fu_370_p2;
wire   [0:0] icmp_ln197_fu_364_p2;
wire   [31:0] s_8_fu_376_p2;
wire  signed [31:0] icmp_ln118_fu_412_p0;
wire  signed [31:0] icmp_ln120_fu_418_p0;
wire  signed [31:0] icmp_ln121_fu_424_p0;
wire  signed [31:0] icmp_ln121_fu_424_p1;
wire   [31:0] select_ln193_1_fu_391_p3;
wire  signed [31:0] sext_ln122_fu_436_p0;
wire  signed [32:0] sext_ln122_fu_436_p1;
wire  signed [31:0] sext_ln122_2_fu_446_p0;
wire  signed [32:0] sext_ln122_2_fu_446_p1;
wire   [32:0] sub_ln122_fu_440_p2;
wire   [31:0] select_ln193_2_fu_398_p3;
wire   [0:0] icmp_ln122_fu_450_p2;
wire   [31:0] add_ln122_fu_456_p2;
wire   [0:0] icmp_ln118_fu_412_p2;
wire   [0:0] icmp_ln120_fu_418_p2;
wire   [0:0] or_ln120_fu_470_p2;
wire   [0:0] icmp_ln121_fu_424_p2;
wire   [0:0] or_ln121_fu_476_p2;
wire   [31:0] n_4_fu_462_p3;
wire   [0:0] xor_ln121_fu_490_p2;
wire   [0:0] or_ln121_2_fu_496_p2;
wire   [31:0] p_5_fu_430_p2;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ready_sig;
wire    ap_done_sig;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 n_3_fu_66 = 32'd0;
#0 p_fu_70 = 32'd0;
#0 c_fu_74 = 31'd0;
#0 s_5_fu_78 = 32'd0;
#0 j_fu_82 = 64'd0;
#0 indvar_flatten8_fu_86 = 95'd0;
#0 ap_done_reg = 1'b0;
end

fmm_reduce_kernel_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready_sig),
    .ap_done(ap_done_sig),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b0 == ap_block_pp0_stage0_subdone) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter2_reg == 1'b0))) begin
        ap_loop_exit_ready_pp0_iter3_reg <= 1'b0;
    end else if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            c_fu_74 <= 31'd0;
        end else if (((icmp_ln192_fu_201_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            c_fu_74 <= add_ln115_fu_249_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            indvar_flatten8_fu_86 <= 95'd0;
        end else if (((icmp_ln192_fu_201_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            indvar_flatten8_fu_86 <= add_ln192_fu_206_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        if ((ap_loop_init == 1'b1)) begin
            j_fu_82 <= zext_ln192_cast_fu_152_p1;
        end else if (((icmp_ln192_fu_201_p2 == 1'd0) & (ap_enable_reg_pp0_iter1 == 1'b1))) begin
            j_fu_82 <= select_ln192_fu_229_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            n_3_fu_66 <= 32'd0;
        end else if (((icmp_ln192_reg_589_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
            n_3_fu_66 <= n_5_fu_482_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            p_fu_70 <= 32'd0;
        end else if (((icmp_ln192_reg_589_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
            p_fu_70 <= p_6_fu_502_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        if (((1'b1 == ap_CS_fsm_pp0_stage0) & (ap_loop_init == 1'b1))) begin
            s_5_fu_78 <= s_4;
        end else if (((icmp_ln192_reg_589_pp0_iter2_reg == 1'd0) & (ap_enable_reg_pp0_iter3 == 1'b1))) begin
            s_5_fu_78 <= select_ln192_1_fu_405_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        icmp_ln115_reg_582 <= icmp_ln115_fu_196_p2;
        icmp_ln192_reg_589 <= icmp_ln192_fu_201_p2;
        trunc_ln117_reg_603 <= trunc_ln117_fu_245_p1;
        trunc_ln119_2_reg_598 <= trunc_ln119_2_fu_241_p1;
        trunc_ln119_reg_593 <= trunc_ln119_fu_237_p1;
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        icmp_ln115_reg_582_pp0_iter2_reg <= icmp_ln115_reg_582;
        icmp_ln192_reg_589_pp0_iter2_reg <= icmp_ln192_reg_589;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        M_e_ce0_local = 1'b1;
    end else begin
        M_e_ce0_local = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_11001) & (ap_enable_reg_pp0_iter2 == 1'b1))) begin
        M_e_ce1_local = 1'b1;
    end else begin
        M_e_ce1_local = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln192_fu_201_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_start_int == 1'b0) & (ap_idle_pp0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((1'b0 == ap_block_pp0_stage0_subdone) & (ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln192_reg_589_pp0_iter2_reg == 1'd1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_loop_exit_ready_pp0_iter3_reg == 1'b1))) begin
        s_9_out_ap_vld = 1'b1;
    end else begin
        s_9_out_ap_vld = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign M_e_address0 = zext_ln119_fu_304_p1;

assign M_e_address1 = zext_ln117_fu_294_p1;

assign M_e_ce0 = M_e_ce0_local;

assign M_e_ce1 = M_e_ce1_local;

assign add_ln115_fu_249_p2 = (select_ln193_fu_221_p3 + 31'd1);

assign add_ln117_fu_290_p2 = (mul_ln117_1 + trunc_ln117_reg_603);

assign add_ln119_2_fu_299_p2 = (add_ln119_fu_284_p2 + trunc_ln117_reg_603);

assign add_ln119_fu_284_p2 = (p_shl_fu_270_p3 + p_shl4_fu_277_p3);

assign add_ln122_fu_456_p2 = (select_ln193_2_fu_398_p3 + 32'd1);

assign add_ln192_1_fu_215_p2 = (j_fu_82 + 64'd1);

assign add_ln192_fu_206_p2 = (indvar_flatten8_fu_86 + 95'd1);

assign add_ln196_fu_334_p2 = ($signed(p_fu_70) + $signed(32'd4294967295));

assign add_ln197_fu_370_p2 = ($signed(s_7_fu_346_p3) + $signed(32'd4294967295));

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_01001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_11001 = ~(1'b1 == 1'b1);

assign ap_block_pp0_stage0_subdone = ~(1'b1 == 1'b1);

assign ap_done = ap_done_sig;

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign ap_ready = ap_ready_sig;

assign icmp_ln115_fu_196_p2 = (($signed(zext_ln115_fu_192_p1) < $signed(cols_non_t)) ? 1'b1 : 1'b0);

assign icmp_ln118_fu_412_p0 = M_e_q1;

assign icmp_ln118_fu_412_p2 = ((icmp_ln118_fu_412_p0 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln120_fu_418_p0 = M_e_q0;

assign icmp_ln120_fu_418_p2 = ((icmp_ln120_fu_418_p0 == 32'd0) ? 1'b1 : 1'b0);

assign icmp_ln121_fu_424_p0 = M_e_q1;

assign icmp_ln121_fu_424_p1 = M_e_q0;

assign icmp_ln121_fu_424_p2 = ((icmp_ln121_fu_424_p0 == icmp_ln121_fu_424_p1) ? 1'b1 : 1'b0);

assign icmp_ln122_fu_450_p2 = ((sext_ln122_2_fu_446_p1 == sub_ln122_fu_440_p2) ? 1'b1 : 1'b0);

assign icmp_ln192_fu_201_p2 = ((indvar_flatten8_fu_86 == mul_ln191) ? 1'b1 : 1'b0);

assign icmp_ln196_fu_328_p2 = (($signed(tmp_fu_318_p4) > $signed(31'd0)) ? 1'b1 : 1'b0);

assign icmp_ln197_fu_364_p2 = (($signed(tmp_3_fu_354_p4) > $signed(31'd0)) ? 1'b1 : 1'b0);

assign n_4_fu_462_p3 = ((icmp_ln122_fu_450_p2[0:0] == 1'b1) ? add_ln122_fu_456_p2 : select_ln193_2_fu_398_p3);

assign n_5_fu_482_p3 = ((or_ln121_fu_476_p2[0:0] == 1'b1) ? select_ln193_2_fu_398_p3 : n_4_fu_462_p3);

assign or_ln120_fu_470_p2 = (icmp_ln120_fu_418_p2 | icmp_ln118_fu_412_p2);

assign or_ln121_2_fu_496_p2 = (xor_ln121_fu_490_p2 | or_ln120_fu_470_p2);

assign or_ln121_fu_476_p2 = (or_ln120_fu_470_p2 | icmp_ln121_fu_424_p2);

assign p_5_fu_430_p2 = (select_ln193_1_fu_391_p3 + 32'd1);

assign p_6_fu_502_p3 = ((or_ln121_2_fu_496_p2[0:0] == 1'b1) ? select_ln193_1_fu_391_p3 : p_5_fu_430_p2);

assign p_shl4_fu_277_p3 = {{trunc_ln119_2_reg_598}, {6'd0}};

assign p_shl_fu_270_p3 = {{trunc_ln119_reg_593}, {8'd0}};

assign s_6_fu_340_p2 = (add_ln196_fu_334_p2 + s_5_fu_78);

assign s_7_fu_346_p3 = ((icmp_ln196_fu_328_p2[0:0] == 1'b1) ? s_6_fu_340_p2 : s_5_fu_78);

assign s_8_fu_376_p2 = (add_ln197_fu_370_p2 + n_3_fu_66);

assign s_9_fu_382_p3 = ((icmp_ln197_fu_364_p2[0:0] == 1'b1) ? s_8_fu_376_p2 : s_7_fu_346_p3);

assign s_9_out = s_9_fu_382_p3;

assign select_ln192_1_fu_405_p3 = ((icmp_ln115_reg_582_pp0_iter2_reg[0:0] == 1'b1) ? s_5_fu_78 : s_9_fu_382_p3);

assign select_ln192_fu_229_p3 = ((icmp_ln115_fu_196_p2[0:0] == 1'b1) ? j_fu_82 : add_ln192_1_fu_215_p2);

assign select_ln193_1_fu_391_p3 = ((icmp_ln115_reg_582_pp0_iter2_reg[0:0] == 1'b1) ? p_fu_70 : 32'd0);

assign select_ln193_2_fu_398_p3 = ((icmp_ln115_reg_582_pp0_iter2_reg[0:0] == 1'b1) ? n_3_fu_66 : 32'd0);

assign select_ln193_fu_221_p3 = ((icmp_ln115_fu_196_p2[0:0] == 1'b1) ? c_fu_74 : 31'd0);

assign sext_ln122_2_fu_446_p0 = M_e_q1;

assign sext_ln122_2_fu_446_p1 = sext_ln122_2_fu_446_p0;

assign sext_ln122_fu_436_p0 = M_e_q0;

assign sext_ln122_fu_436_p1 = sext_ln122_fu_436_p0;

assign sub_ln122_fu_440_p2 = ($signed(33'd0) - $signed(sext_ln122_fu_436_p1));

assign tmp_3_fu_354_p4 = {{n_3_fu_66[31:1]}};

assign tmp_fu_318_p4 = {{p_fu_70[31:1]}};

assign trunc_ln117_fu_245_p1 = select_ln193_fu_221_p3[16:0];

assign trunc_ln119_2_fu_241_p1 = select_ln192_fu_229_p3[10:0];

assign trunc_ln119_fu_237_p1 = select_ln192_fu_229_p3[8:0];

assign xor_ln121_fu_490_p2 = (icmp_ln121_fu_424_p2 ^ 1'd1);

assign zext_ln115_fu_192_p1 = c_fu_74;

assign zext_ln117_fu_294_p1 = add_ln117_fu_290_p2;

assign zext_ln119_fu_304_p1 = add_ln119_2_fu_299_p2;

assign zext_ln192_cast_fu_152_p1 = zext_ln192;

endmodule //fmm_reduce_kernel_greedy_potential_reduce_with_debug_Pipeline_VITIS_LOOP_192_2_VITIS_LOOP_115_1
