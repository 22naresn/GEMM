`timescale 1 ns / 1 ps 

module fmm_reduce_kernel_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4 (
        ap_clk,
        ap_rst,
        ap_start,
        ap_done,
        ap_idle,
        ap_ready,
        m_axi_gmem_0_AWVALID,
        m_axi_gmem_0_AWREADY,
        m_axi_gmem_0_AWADDR,
        m_axi_gmem_0_AWID,
        m_axi_gmem_0_AWLEN,
        m_axi_gmem_0_AWSIZE,
        m_axi_gmem_0_AWBURST,
        m_axi_gmem_0_AWLOCK,
        m_axi_gmem_0_AWCACHE,
        m_axi_gmem_0_AWPROT,
        m_axi_gmem_0_AWQOS,
        m_axi_gmem_0_AWREGION,
        m_axi_gmem_0_AWUSER,
        m_axi_gmem_0_WVALID,
        m_axi_gmem_0_WREADY,
        m_axi_gmem_0_WDATA,
        m_axi_gmem_0_WSTRB,
        m_axi_gmem_0_WLAST,
        m_axi_gmem_0_WID,
        m_axi_gmem_0_WUSER,
        m_axi_gmem_0_ARVALID,
        m_axi_gmem_0_ARREADY,
        m_axi_gmem_0_ARADDR,
        m_axi_gmem_0_ARID,
        m_axi_gmem_0_ARLEN,
        m_axi_gmem_0_ARSIZE,
        m_axi_gmem_0_ARBURST,
        m_axi_gmem_0_ARLOCK,
        m_axi_gmem_0_ARCACHE,
        m_axi_gmem_0_ARPROT,
        m_axi_gmem_0_ARQOS,
        m_axi_gmem_0_ARREGION,
        m_axi_gmem_0_ARUSER,
        m_axi_gmem_0_RVALID,
        m_axi_gmem_0_RREADY,
        m_axi_gmem_0_RDATA,
        m_axi_gmem_0_RLAST,
        m_axi_gmem_0_RID,
        m_axi_gmem_0_RFIFONUM,
        m_axi_gmem_0_RUSER,
        m_axi_gmem_0_RRESP,
        m_axi_gmem_0_BVALID,
        m_axi_gmem_0_BREADY,
        m_axi_gmem_0_BRESP,
        m_axi_gmem_0_BID,
        m_axi_gmem_0_BUSER,
        cols,
        mul_ln58,
        A_dram,
        sext_ln58,
        M_e_address0,
        M_e_ce0,
        M_e_we0,
        M_e_d0
);

parameter    ap_ST_fsm_pp0_stage0 = 1'd1;

input   ap_clk;
input   ap_rst;
input   ap_start;
output   ap_done;
output   ap_idle;
output   ap_ready;
output   m_axi_gmem_0_AWVALID;
input   m_axi_gmem_0_AWREADY;
output  [63:0] m_axi_gmem_0_AWADDR;
output  [0:0] m_axi_gmem_0_AWID;
output  [31:0] m_axi_gmem_0_AWLEN;
output  [2:0] m_axi_gmem_0_AWSIZE;
output  [1:0] m_axi_gmem_0_AWBURST;
output  [1:0] m_axi_gmem_0_AWLOCK;
output  [3:0] m_axi_gmem_0_AWCACHE;
output  [2:0] m_axi_gmem_0_AWPROT;
output  [3:0] m_axi_gmem_0_AWQOS;
output  [3:0] m_axi_gmem_0_AWREGION;
output  [0:0] m_axi_gmem_0_AWUSER;
output   m_axi_gmem_0_WVALID;
input   m_axi_gmem_0_WREADY;
output  [31:0] m_axi_gmem_0_WDATA;
output  [3:0] m_axi_gmem_0_WSTRB;
output   m_axi_gmem_0_WLAST;
output  [0:0] m_axi_gmem_0_WID;
output  [0:0] m_axi_gmem_0_WUSER;
output   m_axi_gmem_0_ARVALID;
input   m_axi_gmem_0_ARREADY;
output  [63:0] m_axi_gmem_0_ARADDR;
output  [0:0] m_axi_gmem_0_ARID;
output  [31:0] m_axi_gmem_0_ARLEN;
output  [2:0] m_axi_gmem_0_ARSIZE;
output  [1:0] m_axi_gmem_0_ARBURST;
output  [1:0] m_axi_gmem_0_ARLOCK;
output  [3:0] m_axi_gmem_0_ARCACHE;
output  [2:0] m_axi_gmem_0_ARPROT;
output  [3:0] m_axi_gmem_0_ARQOS;
output  [3:0] m_axi_gmem_0_ARREGION;
output  [0:0] m_axi_gmem_0_ARUSER;
input   m_axi_gmem_0_RVALID;
output   m_axi_gmem_0_RREADY;
input  [31:0] m_axi_gmem_0_RDATA;
input   m_axi_gmem_0_RLAST;
input  [0:0] m_axi_gmem_0_RID;
input  [8:0] m_axi_gmem_0_RFIFONUM;
input  [0:0] m_axi_gmem_0_RUSER;
input  [1:0] m_axi_gmem_0_RRESP;
input   m_axi_gmem_0_BVALID;
output   m_axi_gmem_0_BREADY;
input  [1:0] m_axi_gmem_0_BRESP;
input  [0:0] m_axi_gmem_0_BID;
input  [0:0] m_axi_gmem_0_BUSER;
input  [31:0] cols;
input  [61:0] mul_ln58;
input  [63:0] A_dram;
input  [31:0] sext_ln58;
output  [16:0] M_e_address0;
output   M_e_ce0;
output   M_e_we0;
output  [31:0] M_e_d0;

reg ap_idle;
reg m_axi_gmem_0_ARVALID;
reg m_axi_gmem_0_RREADY;

(* fsm_encoding = "none" *) reg   [0:0] ap_CS_fsm;
wire    ap_CS_fsm_pp0_stage0;
wire    ap_enable_reg_pp0_iter0;
reg    ap_enable_reg_pp0_iter1;
reg    ap_enable_reg_pp0_iter2;
reg    ap_enable_reg_pp0_iter3;
reg    ap_enable_reg_pp0_iter4;
reg    ap_enable_reg_pp0_iter5;
reg    ap_enable_reg_pp0_iter6;
reg    ap_enable_reg_pp0_iter7;
reg    ap_enable_reg_pp0_iter8;
reg    ap_enable_reg_pp0_iter9;
reg    ap_enable_reg_pp0_iter10;
reg    ap_enable_reg_pp0_iter11;
reg    ap_enable_reg_pp0_iter12;
reg    ap_enable_reg_pp0_iter13;
reg    ap_idle_pp0;
reg   [0:0] icmp_ln58_reg_400;
reg   [0:0] icmp_ln58_reg_400_pp0_iter3_reg;
reg   [0:0] icmp_ln62_reg_434;
reg    ap_predicate_op68_readreq_state5;
reg    ap_block_state5_io;
reg   [0:0] icmp_ln58_reg_400_pp0_iter11_reg;
reg   [0:0] icmp_ln62_reg_434_pp0_iter11_reg;
reg    ap_predicate_op76_read_state13;
reg    ap_block_state13_pp0_stage0_iter12;
reg    ap_block_pp0_stage0_subdone;
wire   [0:0] icmp_ln58_fu_194_p2;
reg    ap_condition_exit_pp0_iter1_stage0;
wire    ap_loop_exit_ready;
reg    ap_ready_int;
reg    gmem_blk_n_AR;
wire    ap_block_pp0_stage0;
reg    gmem_blk_n_R;
reg    ap_block_pp0_stage0_11001;
wire  signed [61:0] sext_ln58_cast_fu_160_p1;
reg  signed [61:0] sext_ln58_cast_reg_395;
reg   [0:0] icmp_ln58_reg_400_pp0_iter2_reg;
reg   [0:0] icmp_ln58_reg_400_pp0_iter4_reg;
reg   [0:0] icmp_ln58_reg_400_pp0_iter5_reg;
reg   [0:0] icmp_ln58_reg_400_pp0_iter6_reg;
reg   [0:0] icmp_ln58_reg_400_pp0_iter7_reg;
reg   [0:0] icmp_ln58_reg_400_pp0_iter8_reg;
reg   [0:0] icmp_ln58_reg_400_pp0_iter9_reg;
reg   [0:0] icmp_ln58_reg_400_pp0_iter10_reg;
reg   [0:0] icmp_ln58_reg_400_pp0_iter12_reg;
wire   [30:0] select_ln58_fu_214_p3;
reg   [30:0] select_ln58_reg_404;
reg   [30:0] select_ln58_reg_404_pp0_iter2_reg;
wire   [30:0] select_ln58_1_fu_222_p3;
reg   [30:0] select_ln58_1_reg_409;
wire   [16:0] trunc_ln65_2_fu_260_p1;
reg   [16:0] trunc_ln65_2_reg_414;
wire   [16:0] trunc_ln65_3_fu_264_p1;
reg   [16:0] trunc_ln65_3_reg_419;
wire   [61:0] empty_fu_156_p2;
reg   [61:0] empty_reg_424;
reg   [16:0] M_e_addr_reg_429;
reg   [16:0] M_e_addr_reg_429_pp0_iter3_reg;
reg   [16:0] M_e_addr_reg_429_pp0_iter4_reg;
reg   [16:0] M_e_addr_reg_429_pp0_iter5_reg;
reg   [16:0] M_e_addr_reg_429_pp0_iter6_reg;
reg   [16:0] M_e_addr_reg_429_pp0_iter7_reg;
reg   [16:0] M_e_addr_reg_429_pp0_iter8_reg;
reg   [16:0] M_e_addr_reg_429_pp0_iter9_reg;
reg   [16:0] M_e_addr_reg_429_pp0_iter10_reg;
reg   [16:0] M_e_addr_reg_429_pp0_iter11_reg;
reg   [16:0] M_e_addr_reg_429_pp0_iter12_reg;
wire   [0:0] icmp_ln62_fu_320_p2;
reg   [0:0] icmp_ln62_reg_434_pp0_iter4_reg;
reg   [0:0] icmp_ln62_reg_434_pp0_iter5_reg;
reg   [0:0] icmp_ln62_reg_434_pp0_iter6_reg;
reg   [0:0] icmp_ln62_reg_434_pp0_iter7_reg;
reg   [0:0] icmp_ln62_reg_434_pp0_iter8_reg;
reg   [0:0] icmp_ln62_reg_434_pp0_iter9_reg;
reg   [0:0] icmp_ln62_reg_434_pp0_iter10_reg;
reg   [0:0] icmp_ln62_reg_434_pp0_iter12_reg;
reg   [63:0] gmem_addr_reg_438;
reg   [31:0] gmem_addr_read_reg_444;
reg   [31:0] ap_phi_mux_storemerge_i_phi_fu_148_p4;
reg   [31:0] ap_phi_reg_pp0_iter13_storemerge_i_reg_144;
wire   [31:0] ap_phi_reg_pp0_iter0_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter1_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter2_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter3_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter4_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter5_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter6_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter7_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter8_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter9_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter10_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter11_storemerge_i_reg_144;
reg   [31:0] ap_phi_reg_pp0_iter12_storemerge_i_reg_144;
wire   [63:0] zext_ln65_fu_297_p1;
wire  signed [63:0] sext_ln63_fu_349_p1;
reg   [30:0] c_1_fu_84;
wire   [30:0] add_ln59_fu_268_p2;
wire    ap_loop_init;
reg   [30:0] r_fu_88;
reg   [61:0] indvar_flatten7_fu_92;
wire   [61:0] add_ln58_1_fu_199_p2;
reg    M_e_we0_local;
reg    M_e_ce0_local;
wire  signed [31:0] empty_fu_156_p0;
wire   [30:0] empty_fu_156_p1;
wire   [31:0] zext_ln59_fu_185_p1;
wire   [0:0] icmp_ln59_fu_189_p2;
wire   [30:0] add_ln58_fu_208_p2;
wire   [26:0] trunc_ln65_fu_230_p1;
wire   [28:0] trunc_ln65_1_fu_242_p1;
wire   [34:0] p_shl_fu_234_p3;
wire   [34:0] p_shl2_fu_246_p3;
wire   [34:0] add_ln65_1_fu_254_p2;
wire   [16:0] add_ln65_fu_293_p2;
wire   [61:0] zext_ln59_1_fu_302_p1;
wire   [61:0] add_ln61_fu_305_p2;
wire   [15:0] tmp_fu_310_p4;
wire   [63:0] shl_ln_fu_326_p3;
wire   [63:0] add_ln63_fu_334_p2;
wire   [61:0] trunc_ln2_fu_339_p4;
reg    ap_done_reg;
wire    ap_continue_int;
reg    ap_done_int;
reg    ap_loop_exit_ready_pp0_iter2_reg;
reg    ap_loop_exit_ready_pp0_iter3_reg;
reg    ap_loop_exit_ready_pp0_iter4_reg;
reg    ap_loop_exit_ready_pp0_iter5_reg;
reg    ap_loop_exit_ready_pp0_iter6_reg;
reg    ap_loop_exit_ready_pp0_iter7_reg;
reg    ap_loop_exit_ready_pp0_iter8_reg;
reg    ap_loop_exit_ready_pp0_iter9_reg;
reg    ap_loop_exit_ready_pp0_iter10_reg;
reg    ap_loop_exit_ready_pp0_iter11_reg;
reg    ap_loop_exit_ready_pp0_iter12_reg;
reg   [0:0] ap_NS_fsm;
wire    ap_enable_pp0;
wire    ap_start_int;
wire    ap_ready_sig;
wire    ap_done_sig;
wire   [61:0] empty_fu_156_p10;
wire    ap_ce_reg;

// power-on initialization
initial begin
#0 ap_CS_fsm = 1'd1;
#0 ap_enable_reg_pp0_iter1 = 1'b0;
#0 ap_enable_reg_pp0_iter2 = 1'b0;
#0 ap_enable_reg_pp0_iter3 = 1'b0;
#0 ap_enable_reg_pp0_iter4 = 1'b0;
#0 ap_enable_reg_pp0_iter5 = 1'b0;
#0 ap_enable_reg_pp0_iter6 = 1'b0;
#0 ap_enable_reg_pp0_iter7 = 1'b0;
#0 ap_enable_reg_pp0_iter8 = 1'b0;
#0 ap_enable_reg_pp0_iter9 = 1'b0;
#0 ap_enable_reg_pp0_iter10 = 1'b0;
#0 ap_enable_reg_pp0_iter11 = 1'b0;
#0 ap_enable_reg_pp0_iter12 = 1'b0;
#0 ap_enable_reg_pp0_iter13 = 1'b0;
#0 c_1_fu_84 = 31'd0;
#0 r_fu_88 = 31'd0;
#0 indvar_flatten7_fu_92 = 62'd0;
#0 ap_done_reg = 1'b0;
end

fmm_reduce_kernel_mul_32s_31ns_62_1_1 #(
    .ID( 1 ),
    .NUM_STAGE( 1 ),
    .din0_WIDTH( 32 ),
    .din1_WIDTH( 31 ),
    .dout_WIDTH( 62 ))
mul_32s_31ns_62_1_1_U20(
    .din0(empty_fu_156_p0),
    .din1(empty_fu_156_p1),
    .dout(empty_fu_156_p2)
);

fmm_reduce_kernel_flow_control_loop_pipe_sequential_init flow_control_loop_pipe_sequential_init_U(
    .ap_clk(ap_clk),
    .ap_rst(ap_rst),
    .ap_start(ap_start),
    .ap_ready(ap_ready_sig),
    .ap_done(ap_done_sig),
    .ap_start_int(ap_start_int),
    .ap_loop_init(ap_loop_init),
    .ap_ready_int(ap_ready_int),
    .ap_loop_exit_ready(ap_condition_exit_pp0_iter1_stage0),
    .ap_loop_exit_done(ap_done_int),
    .ap_continue_int(ap_continue_int),
    .ap_done_int(ap_done_int)
);

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_CS_fsm <= ap_ST_fsm_pp0_stage0;
    end else begin
        ap_CS_fsm <= ap_NS_fsm;
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_done_reg <= 1'b0;
    end else begin
        if ((ap_continue_int == 1'b1)) begin
            ap_done_reg <= 1'b0;
        end else if (((ap_loop_exit_ready_pp0_iter12_reg == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_done_reg <= 1'b1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter1 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter1 <= 1'b0;
        end else if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
            ap_enable_reg_pp0_iter1 <= ap_start_int;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter10 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter10 <= ap_enable_reg_pp0_iter9;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter11 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter11 <= ap_enable_reg_pp0_iter10;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter12 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter12 <= ap_enable_reg_pp0_iter11;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter13 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter13 <= ap_enable_reg_pp0_iter12;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter2 <= 1'b0;
    end else begin
        if ((1'b1 == ap_condition_exit_pp0_iter1_stage0)) begin
            ap_enable_reg_pp0_iter2 <= 1'b0;
        end else if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter2 <= ap_enable_reg_pp0_iter1;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter3 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter3 <= ap_enable_reg_pp0_iter2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter4 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter4 <= ap_enable_reg_pp0_iter3;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter5 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter5 <= ap_enable_reg_pp0_iter4;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter6 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter6 <= ap_enable_reg_pp0_iter5;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter7 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter7 <= ap_enable_reg_pp0_iter6;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter8 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter8 <= ap_enable_reg_pp0_iter7;
        end
    end
end

always @ (posedge ap_clk) begin
    if (ap_rst == 1'b1) begin
        ap_enable_reg_pp0_iter9 <= 1'b0;
    end else begin
        if ((1'b0 == ap_block_pp0_stage0_subdone)) begin
            ap_enable_reg_pp0_iter9 <= ap_enable_reg_pp0_iter8;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter3 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        if (((icmp_ln62_fu_320_p2 == 1'd0) & (icmp_ln58_reg_400_pp0_iter2_reg == 1'd0))) begin
            ap_phi_reg_pp0_iter4_storemerge_i_reg_144 <= 32'd0;
        end else if ((1'b1 == 1'b1)) begin
            ap_phi_reg_pp0_iter4_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter3_storemerge_i_reg_144;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        if ((ap_loop_init == 1'b1)) begin
            c_1_fu_84 <= 31'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln58_fu_194_p2 == 1'd0))) begin
            c_1_fu_84 <= add_ln59_fu_268_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        if ((ap_loop_init == 1'b1)) begin
            indvar_flatten7_fu_92 <= 62'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln58_fu_194_p2 == 1'd0))) begin
            indvar_flatten7_fu_92 <= add_ln58_1_fu_199_p2;
        end
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        if ((ap_loop_init == 1'b1)) begin
            r_fu_88 <= 31'd0;
        end else if (((ap_enable_reg_pp0_iter1 == 1'b1) & (icmp_ln58_fu_194_p2 == 1'd0))) begin
            r_fu_88 <= select_ln58_1_fu_222_p3;
        end
    end
end

always @ (posedge ap_clk) begin
    if ((1'b0 == ap_block_pp0_stage0_11001)) begin
        M_e_addr_reg_429 <= zext_ln65_fu_297_p1;
        M_e_addr_reg_429_pp0_iter10_reg <= M_e_addr_reg_429_pp0_iter9_reg;
        M_e_addr_reg_429_pp0_iter11_reg <= M_e_addr_reg_429_pp0_iter10_reg;
        M_e_addr_reg_429_pp0_iter12_reg <= M_e_addr_reg_429_pp0_iter11_reg;
        M_e_addr_reg_429_pp0_iter3_reg <= M_e_addr_reg_429;
        M_e_addr_reg_429_pp0_iter4_reg <= M_e_addr_reg_429_pp0_iter3_reg;
        M_e_addr_reg_429_pp0_iter5_reg <= M_e_addr_reg_429_pp0_iter4_reg;
        M_e_addr_reg_429_pp0_iter6_reg <= M_e_addr_reg_429_pp0_iter5_reg;
        M_e_addr_reg_429_pp0_iter7_reg <= M_e_addr_reg_429_pp0_iter6_reg;
        M_e_addr_reg_429_pp0_iter8_reg <= M_e_addr_reg_429_pp0_iter7_reg;
        M_e_addr_reg_429_pp0_iter9_reg <= M_e_addr_reg_429_pp0_iter8_reg;
        ap_loop_exit_ready_pp0_iter10_reg <= ap_loop_exit_ready_pp0_iter9_reg;
        ap_loop_exit_ready_pp0_iter11_reg <= ap_loop_exit_ready_pp0_iter10_reg;
        ap_loop_exit_ready_pp0_iter12_reg <= ap_loop_exit_ready_pp0_iter11_reg;
        ap_loop_exit_ready_pp0_iter3_reg <= ap_loop_exit_ready_pp0_iter2_reg;
        ap_loop_exit_ready_pp0_iter4_reg <= ap_loop_exit_ready_pp0_iter3_reg;
        ap_loop_exit_ready_pp0_iter5_reg <= ap_loop_exit_ready_pp0_iter4_reg;
        ap_loop_exit_ready_pp0_iter6_reg <= ap_loop_exit_ready_pp0_iter5_reg;
        ap_loop_exit_ready_pp0_iter7_reg <= ap_loop_exit_ready_pp0_iter6_reg;
        ap_loop_exit_ready_pp0_iter8_reg <= ap_loop_exit_ready_pp0_iter7_reg;
        ap_loop_exit_ready_pp0_iter9_reg <= ap_loop_exit_ready_pp0_iter8_reg;
        empty_reg_424 <= empty_fu_156_p2;
        gmem_addr_read_reg_444 <= m_axi_gmem_0_RDATA;
        gmem_addr_reg_438 <= sext_ln63_fu_349_p1;
        icmp_ln58_reg_400_pp0_iter10_reg <= icmp_ln58_reg_400_pp0_iter9_reg;
        icmp_ln58_reg_400_pp0_iter11_reg <= icmp_ln58_reg_400_pp0_iter10_reg;
        icmp_ln58_reg_400_pp0_iter12_reg <= icmp_ln58_reg_400_pp0_iter11_reg;
        icmp_ln58_reg_400_pp0_iter2_reg <= icmp_ln58_reg_400;
        icmp_ln58_reg_400_pp0_iter3_reg <= icmp_ln58_reg_400_pp0_iter2_reg;
        icmp_ln58_reg_400_pp0_iter4_reg <= icmp_ln58_reg_400_pp0_iter3_reg;
        icmp_ln58_reg_400_pp0_iter5_reg <= icmp_ln58_reg_400_pp0_iter4_reg;
        icmp_ln58_reg_400_pp0_iter6_reg <= icmp_ln58_reg_400_pp0_iter5_reg;
        icmp_ln58_reg_400_pp0_iter7_reg <= icmp_ln58_reg_400_pp0_iter6_reg;
        icmp_ln58_reg_400_pp0_iter8_reg <= icmp_ln58_reg_400_pp0_iter7_reg;
        icmp_ln58_reg_400_pp0_iter9_reg <= icmp_ln58_reg_400_pp0_iter8_reg;
        icmp_ln62_reg_434 <= icmp_ln62_fu_320_p2;
        icmp_ln62_reg_434_pp0_iter10_reg <= icmp_ln62_reg_434_pp0_iter9_reg;
        icmp_ln62_reg_434_pp0_iter11_reg <= icmp_ln62_reg_434_pp0_iter10_reg;
        icmp_ln62_reg_434_pp0_iter12_reg <= icmp_ln62_reg_434_pp0_iter11_reg;
        icmp_ln62_reg_434_pp0_iter4_reg <= icmp_ln62_reg_434;
        icmp_ln62_reg_434_pp0_iter5_reg <= icmp_ln62_reg_434_pp0_iter4_reg;
        icmp_ln62_reg_434_pp0_iter6_reg <= icmp_ln62_reg_434_pp0_iter5_reg;
        icmp_ln62_reg_434_pp0_iter7_reg <= icmp_ln62_reg_434_pp0_iter6_reg;
        icmp_ln62_reg_434_pp0_iter8_reg <= icmp_ln62_reg_434_pp0_iter7_reg;
        icmp_ln62_reg_434_pp0_iter9_reg <= icmp_ln62_reg_434_pp0_iter8_reg;
        select_ln58_reg_404_pp0_iter2_reg <= select_ln58_reg_404;
    end
end

always @ (posedge ap_clk) begin
    if (((1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_loop_exit_ready_pp0_iter2_reg <= ap_loop_exit_ready;
        icmp_ln58_reg_400 <= icmp_ln58_fu_194_p2;
        select_ln58_1_reg_409 <= select_ln58_1_fu_222_p3;
        select_ln58_reg_404 <= select_ln58_fu_214_p3;
        sext_ln58_cast_reg_395 <= sext_ln58_cast_fu_160_p1;
        trunc_ln65_2_reg_414[16 : 6] <= trunc_ln65_2_fu_260_p1[16 : 6];
        trunc_ln65_3_reg_419 <= trunc_ln65_3_fu_264_p1;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter9 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter10_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter9_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter10 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter11_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter10_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter11 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter12_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter11_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter13_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter12_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter1_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter0_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter2_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter1_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter2 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter3_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter2_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter5_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter4_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter5 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter6_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter5_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter6 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter7_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter6_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter7 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter8_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter7_storemerge_i_reg_144;
    end
end

always @ (posedge ap_clk) begin
    if (((ap_enable_reg_pp0_iter8 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        ap_phi_reg_pp0_iter9_storemerge_i_reg_144 <= ap_phi_reg_pp0_iter8_storemerge_i_reg_144;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        M_e_ce0_local = 1'b1;
    end else begin
        M_e_ce0_local = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001))) begin
        M_e_we0_local = 1'b1;
    end else begin
        M_e_we0_local = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter1 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (icmp_ln58_fu_194_p2 == 1'd1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b1;
    end else begin
        ap_condition_exit_pp0_iter1_stage0 = 1'b0;
    end
end

always @ (*) begin
    if (((ap_loop_exit_ready_pp0_iter12_reg == 1'b1) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_done_int = 1'b1;
    end else begin
        ap_done_int = ap_done_reg;
    end
end

always @ (*) begin
    if (((ap_idle_pp0 == 1'b1) & (ap_start_int == 1'b0) & (1'b1 == ap_CS_fsm_pp0_stage0))) begin
        ap_idle = 1'b1;
    end else begin
        ap_idle = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter13 == 1'b0) & (ap_enable_reg_pp0_iter12 == 1'b0) & (ap_enable_reg_pp0_iter11 == 1'b0) & (ap_enable_reg_pp0_iter10 == 1'b0) & (ap_enable_reg_pp0_iter9 == 1'b0) & (ap_enable_reg_pp0_iter8 == 1'b0) & (ap_enable_reg_pp0_iter7 == 1'b0) & (ap_enable_reg_pp0_iter6 == 1'b0) & (ap_enable_reg_pp0_iter5 == 1'b0) & (ap_enable_reg_pp0_iter4 == 1'b0) & (ap_enable_reg_pp0_iter3 == 1'b0) & (ap_enable_reg_pp0_iter2 == 1'b0) & (ap_enable_reg_pp0_iter1 == 1'b0) & (ap_enable_reg_pp0_iter0 == 1'b0))) begin
        ap_idle_pp0 = 1'b1;
    end else begin
        ap_idle_pp0 = 1'b0;
    end
end

always @ (*) begin
    if (((icmp_ln62_reg_434_pp0_iter12_reg == 1'd1) & (icmp_ln58_reg_400_pp0_iter12_reg == 1'd0))) begin
        ap_phi_mux_storemerge_i_phi_fu_148_p4 = gmem_addr_read_reg_444;
    end else begin
        ap_phi_mux_storemerge_i_phi_fu_148_p4 = ap_phi_reg_pp0_iter13_storemerge_i_reg_144;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter0 == 1'b1) & (1'b1 == ap_CS_fsm_pp0_stage0) & (1'b0 == ap_block_pp0_stage0_subdone))) begin
        ap_ready_int = 1'b1;
    end else begin
        ap_ready_int = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (ap_predicate_op68_readreq_state5 == 1'b1))) begin
        gmem_blk_n_AR = m_axi_gmem_0_ARREADY;
    end else begin
        gmem_blk_n_AR = 1'b1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0) & (ap_predicate_op76_read_state13 == 1'b1))) begin
        gmem_blk_n_R = m_axi_gmem_0_RVALID;
    end else begin
        gmem_blk_n_R = 1'b1;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_predicate_op68_readreq_state5 == 1'b1))) begin
        m_axi_gmem_0_ARVALID = 1'b1;
    end else begin
        m_axi_gmem_0_ARVALID = 1'b0;
    end
end

always @ (*) begin
    if (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b0 == ap_block_pp0_stage0_11001) & (ap_predicate_op76_read_state13 == 1'b1))) begin
        m_axi_gmem_0_RREADY = 1'b1;
    end else begin
        m_axi_gmem_0_RREADY = 1'b0;
    end
end

always @ (*) begin
    case (ap_CS_fsm)
        ap_ST_fsm_pp0_stage0 : begin
            ap_NS_fsm = ap_ST_fsm_pp0_stage0;
        end
        default : begin
            ap_NS_fsm = 'bx;
        end
    endcase
end

assign M_e_address0 = M_e_addr_reg_429_pp0_iter12_reg;

assign M_e_ce0 = M_e_ce0_local;

assign M_e_d0 = ap_phi_mux_storemerge_i_phi_fu_148_p4;

assign M_e_we0 = M_e_we0_local;

assign add_ln58_1_fu_199_p2 = (indvar_flatten7_fu_92 + 62'd1);

assign add_ln58_fu_208_p2 = (r_fu_88 + 31'd1);

assign add_ln59_fu_268_p2 = (select_ln58_fu_214_p3 + 31'd1);

assign add_ln61_fu_305_p2 = (empty_reg_424 + zext_ln59_1_fu_302_p1);

assign add_ln63_fu_334_p2 = (shl_ln_fu_326_p3 + A_dram);

assign add_ln65_1_fu_254_p2 = (p_shl_fu_234_p3 + p_shl2_fu_246_p3);

assign add_ln65_fu_293_p2 = (trunc_ln65_2_reg_414 + trunc_ln65_3_reg_419);

assign ap_CS_fsm_pp0_stage0 = ap_CS_fsm[32'd0];

assign ap_block_pp0_stage0 = ~(1'b1 == 1'b1);

always @ (*) begin
    ap_block_pp0_stage0_11001 = (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b1 == ap_block_state13_pp0_stage0_iter12)) | ((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_block_state5_io)));
end

always @ (*) begin
    ap_block_pp0_stage0_subdone = (((ap_enable_reg_pp0_iter12 == 1'b1) & (1'b1 == ap_block_state13_pp0_stage0_iter12)) | ((ap_enable_reg_pp0_iter4 == 1'b1) & (1'b1 == ap_block_state5_io)));
end

always @ (*) begin
    ap_block_state13_pp0_stage0_iter12 = ((ap_predicate_op76_read_state13 == 1'b1) & (m_axi_gmem_0_RVALID == 1'b0));
end

always @ (*) begin
    ap_block_state5_io = ((m_axi_gmem_0_ARREADY == 1'b0) & (ap_predicate_op68_readreq_state5 == 1'b1));
end

assign ap_done = ap_done_sig;

assign ap_enable_pp0 = (ap_idle_pp0 ^ 1'b1);

assign ap_enable_reg_pp0_iter0 = ap_start_int;

assign ap_loop_exit_ready = ap_condition_exit_pp0_iter1_stage0;

assign ap_phi_reg_pp0_iter0_storemerge_i_reg_144 = 'bx;

always @ (*) begin
    ap_predicate_op68_readreq_state5 = ((icmp_ln62_reg_434 == 1'd1) & (icmp_ln58_reg_400_pp0_iter3_reg == 1'd0));
end

always @ (*) begin
    ap_predicate_op76_read_state13 = ((icmp_ln62_reg_434_pp0_iter11_reg == 1'd1) & (icmp_ln58_reg_400_pp0_iter11_reg == 1'd0));
end

assign ap_ready = ap_ready_sig;

assign empty_fu_156_p0 = sext_ln58_cast_reg_395;

assign empty_fu_156_p1 = empty_fu_156_p10;

assign empty_fu_156_p10 = select_ln58_1_reg_409;

assign icmp_ln58_fu_194_p2 = ((indvar_flatten7_fu_92 == mul_ln58) ? 1'b1 : 1'b0);

assign icmp_ln59_fu_189_p2 = (($signed(zext_ln59_fu_185_p1) < $signed(cols)) ? 1'b1 : 1'b0);

assign icmp_ln62_fu_320_p2 = ((tmp_fu_310_p4 == 16'd0) ? 1'b1 : 1'b0);

assign m_axi_gmem_0_ARADDR = gmem_addr_reg_438;

assign m_axi_gmem_0_ARBURST = 2'd0;

assign m_axi_gmem_0_ARCACHE = 4'd0;

assign m_axi_gmem_0_ARID = 1'd0;

assign m_axi_gmem_0_ARLEN = 64'd1;

assign m_axi_gmem_0_ARLOCK = 2'd0;

assign m_axi_gmem_0_ARPROT = 3'd0;

assign m_axi_gmem_0_ARQOS = 4'd0;

assign m_axi_gmem_0_ARREGION = 4'd0;

assign m_axi_gmem_0_ARSIZE = 3'd0;

assign m_axi_gmem_0_ARUSER = 1'd0;

assign m_axi_gmem_0_AWADDR = 64'd0;

assign m_axi_gmem_0_AWBURST = 2'd0;

assign m_axi_gmem_0_AWCACHE = 4'd0;

assign m_axi_gmem_0_AWID = 1'd0;

assign m_axi_gmem_0_AWLEN = 32'd0;

assign m_axi_gmem_0_AWLOCK = 2'd0;

assign m_axi_gmem_0_AWPROT = 3'd0;

assign m_axi_gmem_0_AWQOS = 4'd0;

assign m_axi_gmem_0_AWREGION = 4'd0;

assign m_axi_gmem_0_AWSIZE = 3'd0;

assign m_axi_gmem_0_AWUSER = 1'd0;

assign m_axi_gmem_0_AWVALID = 1'b0;

assign m_axi_gmem_0_BREADY = 1'b0;

assign m_axi_gmem_0_WDATA = 32'd0;

assign m_axi_gmem_0_WID = 1'd0;

assign m_axi_gmem_0_WLAST = 1'b0;

assign m_axi_gmem_0_WSTRB = 4'd0;

assign m_axi_gmem_0_WUSER = 1'd0;

assign m_axi_gmem_0_WVALID = 1'b0;

assign p_shl2_fu_246_p3 = {{trunc_ln65_1_fu_242_p1}, {6'd0}};

assign p_shl_fu_234_p3 = {{trunc_ln65_fu_230_p1}, {8'd0}};

assign select_ln58_1_fu_222_p3 = ((icmp_ln59_fu_189_p2[0:0] == 1'b1) ? r_fu_88 : add_ln58_fu_208_p2);

assign select_ln58_fu_214_p3 = ((icmp_ln59_fu_189_p2[0:0] == 1'b1) ? c_1_fu_84 : 31'd0);

assign sext_ln58_cast_fu_160_p1 = $signed(sext_ln58);

assign sext_ln63_fu_349_p1 = $signed(trunc_ln2_fu_339_p4);

assign shl_ln_fu_326_p3 = {{add_ln61_fu_305_p2}, {2'd0}};

assign tmp_fu_310_p4 = {{add_ln61_fu_305_p2[31:16]}};

assign trunc_ln2_fu_339_p4 = {{add_ln63_fu_334_p2[63:2]}};

assign trunc_ln65_1_fu_242_p1 = select_ln58_1_fu_222_p3[28:0];

assign trunc_ln65_2_fu_260_p1 = add_ln65_1_fu_254_p2[16:0];

assign trunc_ln65_3_fu_264_p1 = select_ln58_fu_214_p3[16:0];

assign trunc_ln65_fu_230_p1 = select_ln58_1_fu_222_p3[26:0];

assign zext_ln59_1_fu_302_p1 = select_ln58_reg_404_pp0_iter2_reg;

assign zext_ln59_fu_185_p1 = c_1_fu_84;

assign zext_ln65_fu_297_p1 = add_ln65_fu_293_p2;

always @ (posedge ap_clk) begin
    trunc_ln65_2_reg_414[5:0] <= 6'b000000;
end

endmodule //fmm_reduce_kernel_load_matrix_from_dram_safe_Pipeline_VITIS_LOOP_58_3_VITIS_LOOP_59_4
